
// Dual Port ROM

module dice6_rom
#(parameter DATA_WIDTH=1, parameter ADDR_WIDTH=12)
(
	input [(ADDR_WIDTH-1):0] addr,
	input clk, 
	output reg [(DATA_WIDTH-1):0] q
);

	// Declare the ROM variable
	reg [DATA_WIDTH-1:0] rom[2**ADDR_WIDTH-1:0];

   // value to Draw Dine Face 6
	initial
	begin
     rom[0] = 0;
     rom[1] = 0;
     rom[2] = 0;
     rom[3] = 0;
     rom[4] = 0;
     rom[5] = 0;
     rom[6] = 0;
     rom[7] = 0;
     rom[8] = 0;
     rom[9] = 0;
     rom[10] = 0;
     rom[11] = 0;
     rom[12] = 0;
     rom[13] = 0;
     rom[14] = 0;
     rom[15] = 0;
     rom[16] = 0;
     rom[17] = 0;
     rom[18] = 0;
     rom[19] = 0;
     rom[20] = 0;
     rom[21] = 0;
     rom[22] = 0;
     rom[23] = 0;
     rom[24] = 0;
     rom[25] = 0;
     rom[26] = 0;
     rom[27] = 0;
     rom[28] = 0;
     rom[29] = 0;
     rom[30] = 0;
     rom[31] = 0;
     rom[32] = 0;
     rom[33] = 0;
     rom[34] = 0;
     rom[35] = 0;
     rom[36] = 0;
     rom[37] = 0;
     rom[38] = 0;
     rom[39] = 0;
     rom[40] = 0;
     rom[41] = 0;
     rom[42] = 0;
     rom[43] = 0;
     rom[44] = 0;
     rom[45] = 0;
     rom[46] = 0;
     rom[47] = 0;
     rom[48] = 0;
     rom[49] = 0;
     rom[50] = 0;
     rom[51] = 0;
     rom[52] = 0;
     rom[53] = 0;
     rom[54] = 0;
     rom[55] = 0;
     rom[56] = 0;
     rom[57] = 0;
     rom[58] = 0;
     rom[59] = 0;
     rom[60] = 0;
     rom[61] = 0;
     rom[62] = 0;
     rom[63] = 0;
     rom[64] = 0;
     rom[65] = 0;
     rom[66] = 0;
     rom[67] = 0;
     rom[68] = 0;
     rom[69] = 0;
     rom[70] = 0;
     rom[71] = 0;
     rom[72] = 0;
     rom[73] = 0;
     rom[74] = 0;
     rom[75] = 0;
     rom[76] = 0;
     rom[77] = 0;
     rom[78] = 0;
     rom[79] = 0;
     rom[80] = 0;
     rom[81] = 0;
     rom[82] = 0;
     rom[83] = 0;
     rom[84] = 0;
     rom[85] = 0;
     rom[86] = 0;
     rom[87] = 0;
     rom[88] = 0;
     rom[89] = 0;
     rom[90] = 0;
     rom[91] = 0;
     rom[92] = 0;
     rom[93] = 0;
     rom[94] = 0;
     rom[95] = 0;
     rom[96] = 0;
     rom[97] = 0;
     rom[98] = 0;
     rom[99] = 0;
     rom[100] = 0;
     rom[101] = 0;
     rom[102] = 0;
     rom[103] = 0;
     rom[104] = 0;
     rom[105] = 0;
     rom[106] = 0;
     rom[107] = 0;
     rom[108] = 0;
     rom[109] = 0;
     rom[110] = 0;
     rom[111] = 0;
     rom[112] = 0;
     rom[113] = 0;
     rom[114] = 0;
     rom[115] = 0;
     rom[116] = 0;
     rom[117] = 0;
     rom[118] = 0;
     rom[119] = 0;
     rom[120] = 0;
     rom[121] = 0;
     rom[122] = 0;
     rom[123] = 0;
     rom[124] = 0;
     rom[125] = 0;
     rom[126] = 0;
     rom[127] = 0;
     rom[128] = 0;
     rom[129] = 0;
     rom[130] = 0;
     rom[131] = 0;
     rom[132] = 0;
     rom[133] = 0;
     rom[134] = 0;
     rom[135] = 0;
     rom[136] = 0;
     rom[137] = 0;
     rom[138] = 0;
     rom[139] = 0;
     rom[140] = 0;
     rom[141] = 0;
     rom[142] = 0;
     rom[143] = 0;
     rom[144] = 0;
     rom[145] = 0;
     rom[146] = 0;
     rom[147] = 0;
     rom[148] = 0;
     rom[149] = 0;
     rom[150] = 0;
     rom[151] = 0;
     rom[152] = 0;
     rom[153] = 0;
     rom[154] = 0;
     rom[155] = 0;
     rom[156] = 0;
     rom[157] = 0;
     rom[158] = 0;
     rom[159] = 0;
     rom[160] = 0;
     rom[161] = 0;
     rom[162] = 0;
     rom[163] = 0;
     rom[164] = 0;
     rom[165] = 0;
     rom[166] = 0;
     rom[167] = 0;
     rom[168] = 0;
     rom[169] = 0;
     rom[170] = 0;
     rom[171] = 0;
     rom[172] = 0;
     rom[173] = 0;
     rom[174] = 0;
     rom[175] = 0;
     rom[176] = 0;
     rom[177] = 0;
     rom[178] = 0;
     rom[179] = 0;
     rom[180] = 0;
     rom[181] = 0;
     rom[182] = 0;
     rom[183] = 0;
     rom[184] = 0;
     rom[185] = 0;
     rom[186] = 0;
     rom[187] = 0;
     rom[188] = 0;
     rom[189] = 0;
     rom[190] = 0;
     rom[191] = 0;
     rom[192] = 0;
     rom[193] = 0;
     rom[194] = 0;
     rom[195] = 0;
     rom[196] = 0;
     rom[197] = 0;
     rom[198] = 0;
     rom[199] = 0;
     rom[200] = 0;
     rom[201] = 0;
     rom[202] = 0;
     rom[203] = 0;
     rom[204] = 0;
     rom[205] = 0;
     rom[206] = 0;
     rom[207] = 0;
     rom[208] = 0;
     rom[209] = 0;
     rom[210] = 0;
     rom[211] = 0;
     rom[212] = 0;
     rom[213] = 0;
     rom[214] = 0;
     rom[215] = 0;
     rom[216] = 0;
     rom[217] = 0;
     rom[218] = 0;
     rom[219] = 0;
     rom[220] = 0;
     rom[221] = 0;
     rom[222] = 0;
     rom[223] = 0;
     rom[224] = 0;
     rom[225] = 0;
     rom[226] = 0;
     rom[227] = 0;
     rom[228] = 0;
     rom[229] = 0;
     rom[230] = 0;
     rom[231] = 0;
     rom[232] = 0;
     rom[233] = 0;
     rom[234] = 0;
     rom[235] = 0;
     rom[236] = 0;
     rom[237] = 0;
     rom[238] = 0;
     rom[239] = 0;
     rom[240] = 0;
     rom[241] = 0;
     rom[242] = 0;
     rom[243] = 0;
     rom[244] = 0;
     rom[245] = 0;
     rom[246] = 0;
     rom[247] = 0;
     rom[248] = 0;
     rom[249] = 0;
     rom[250] = 0;
     rom[251] = 0;
     rom[252] = 0;
     rom[253] = 0;
     rom[254] = 0;
     rom[255] = 0;
     rom[256] = 0;
     rom[257] = 0;
     rom[258] = 0;
     rom[259] = 0;
     rom[260] = 0;
     rom[261] = 0;
     rom[262] = 0;
     rom[263] = 0;
     rom[264] = 0;
     rom[265] = 0;
     rom[266] = 0;
     rom[267] = 0;
     rom[268] = 0;
     rom[269] = 0;
     rom[270] = 0;
     rom[271] = 0;
     rom[272] = 0;
     rom[273] = 0;
     rom[274] = 0;
     rom[275] = 0;
     rom[276] = 0;
     rom[277] = 0;
     rom[278] = 0;
     rom[279] = 0;
     rom[280] = 0;
     rom[281] = 0;
     rom[282] = 0;
     rom[283] = 0;
     rom[284] = 0;
     rom[285] = 0;
     rom[286] = 0;
     rom[287] = 0;
     rom[288] = 0;
     rom[289] = 0;
     rom[290] = 0;
     rom[291] = 0;
     rom[292] = 0;
     rom[293] = 0;
     rom[294] = 0;
     rom[295] = 0;
     rom[296] = 0;
     rom[297] = 0;
     rom[298] = 0;
     rom[299] = 0;
     rom[300] = 0;
     rom[301] = 0;
     rom[302] = 0;
     rom[303] = 0;
     rom[304] = 0;
     rom[305] = 0;
     rom[306] = 0;
     rom[307] = 0;
     rom[308] = 0;
     rom[309] = 0;
     rom[310] = 0;
     rom[311] = 0;
     rom[312] = 0;
     rom[313] = 0;
     rom[314] = 0;
     rom[315] = 0;
     rom[316] = 0;
     rom[317] = 0;
     rom[318] = 0;
     rom[319] = 0;
     rom[320] = 0;
     rom[321] = 0;
     rom[322] = 0;
     rom[323] = 0;
     rom[324] = 0;
     rom[325] = 0;
     rom[326] = 0;
     rom[327] = 0;
     rom[328] = 0;
     rom[329] = 0;
     rom[330] = 0;
     rom[331] = 0;
     rom[332] = 0;
     rom[333] = 0;
     rom[334] = 0;
     rom[335] = 0;
     rom[336] = 0;
     rom[337] = 0;
     rom[338] = 0;
     rom[339] = 0;
     rom[340] = 0;
     rom[341] = 0;
     rom[342] = 0;
     rom[343] = 0;
     rom[344] = 0;
     rom[345] = 0;
     rom[346] = 0;
     rom[347] = 0;
     rom[348] = 0;
     rom[349] = 0;
     rom[350] = 0;
     rom[351] = 0;
     rom[352] = 0;
     rom[353] = 0;
     rom[354] = 0;
     rom[355] = 0;
     rom[356] = 0;
     rom[357] = 0;
     rom[358] = 0;
     rom[359] = 0;
     rom[360] = 0;
     rom[361] = 0;
     rom[362] = 0;
     rom[363] = 0;
     rom[364] = 0;
     rom[365] = 0;
     rom[366] = 0;
     rom[367] = 0;
     rom[368] = 0;
     rom[369] = 0;
     rom[370] = 0;
     rom[371] = 0;
     rom[372] = 0;
     rom[373] = 0;
     rom[374] = 0;
     rom[375] = 0;
     rom[376] = 0;
     rom[377] = 0;
     rom[378] = 0;
     rom[379] = 0;
     rom[380] = 0;
     rom[381] = 0;
     rom[382] = 0;
     rom[383] = 0;
     rom[384] = 0;
     rom[385] = 0;
     rom[386] = 0;
     rom[387] = 0;
     rom[388] = 0;
     rom[389] = 0;
     rom[390] = 0;
     rom[391] = 0;
     rom[392] = 0;
     rom[393] = 0;
     rom[394] = 0;
     rom[395] = 1;
     rom[396] = 1;
     rom[397] = 1;
     rom[398] = 1;
     rom[399] = 1;
     rom[400] = 0;
     rom[401] = 0;
     rom[402] = 0;
     rom[403] = 0;
     rom[404] = 0;
     rom[405] = 0;
     rom[406] = 0;
     rom[407] = 0;
     rom[408] = 0;
     rom[409] = 0;
     rom[410] = 0;
     rom[411] = 0;
     rom[412] = 0;
     rom[413] = 1;
     rom[414] = 1;
     rom[415] = 1;
     rom[416] = 1;
     rom[417] = 1;
     rom[418] = 1;
     rom[419] = 0;
     rom[420] = 0;
     rom[421] = 0;
     rom[422] = 0;
     rom[423] = 0;
     rom[424] = 0;
     rom[425] = 0;
     rom[426] = 0;
     rom[427] = 0;
     rom[428] = 0;
     rom[429] = 0;
     rom[430] = 0;
     rom[431] = 0;
     rom[432] = 1;
     rom[433] = 1;
     rom[434] = 1;
     rom[435] = 1;
     rom[436] = 1;
     rom[437] = 0;
     rom[438] = 0;
     rom[439] = 0;
     rom[440] = 0;
     rom[441] = 0;
     rom[442] = 0;
     rom[443] = 0;
     rom[444] = 0;
     rom[445] = 0;
     rom[446] = 0;
     rom[447] = 0;
     rom[448] = 0;
     rom[449] = 0;
     rom[450] = 0;
     rom[451] = 0;
     rom[452] = 0;
     rom[453] = 0;
     rom[454] = 0;
     rom[455] = 0;
     rom[456] = 0;
     rom[457] = 1;
     rom[458] = 1;
     rom[459] = 1;
     rom[460] = 1;
     rom[461] = 1;
     rom[462] = 1;
     rom[463] = 1;
     rom[464] = 1;
     rom[465] = 1;
     rom[466] = 0;
     rom[467] = 0;
     rom[468] = 0;
     rom[469] = 0;
     rom[470] = 0;
     rom[471] = 0;
     rom[472] = 0;
     rom[473] = 0;
     rom[474] = 0;
     rom[475] = 1;
     rom[476] = 1;
     rom[477] = 1;
     rom[478] = 1;
     rom[479] = 1;
     rom[480] = 1;
     rom[481] = 1;
     rom[482] = 1;
     rom[483] = 1;
     rom[484] = 0;
     rom[485] = 0;
     rom[486] = 0;
     rom[487] = 0;
     rom[488] = 0;
     rom[489] = 0;
     rom[490] = 0;
     rom[491] = 0;
     rom[492] = 0;
     rom[493] = 0;
     rom[494] = 1;
     rom[495] = 1;
     rom[496] = 1;
     rom[497] = 1;
     rom[498] = 1;
     rom[499] = 1;
     rom[500] = 1;
     rom[501] = 1;
     rom[502] = 1;
     rom[503] = 0;
     rom[504] = 0;
     rom[505] = 0;
     rom[506] = 0;
     rom[507] = 0;
     rom[508] = 0;
     rom[509] = 0;
     rom[510] = 0;
     rom[511] = 0;
     rom[512] = 0;
     rom[513] = 0;
     rom[514] = 0;
     rom[515] = 0;
     rom[516] = 0;
     rom[517] = 0;
     rom[518] = 0;
     rom[519] = 0;
     rom[520] = 1;
     rom[521] = 1;
     rom[522] = 1;
     rom[523] = 1;
     rom[524] = 1;
     rom[525] = 1;
     rom[526] = 1;
     rom[527] = 1;
     rom[528] = 1;
     rom[529] = 1;
     rom[530] = 1;
     rom[531] = 0;
     rom[532] = 0;
     rom[533] = 0;
     rom[534] = 0;
     rom[535] = 0;
     rom[536] = 0;
     rom[537] = 0;
     rom[538] = 1;
     rom[539] = 1;
     rom[540] = 1;
     rom[541] = 1;
     rom[542] = 1;
     rom[543] = 1;
     rom[544] = 1;
     rom[545] = 1;
     rom[546] = 1;
     rom[547] = 1;
     rom[548] = 1;
     rom[549] = 1;
     rom[550] = 0;
     rom[551] = 0;
     rom[552] = 0;
     rom[553] = 0;
     rom[554] = 0;
     rom[555] = 0;
     rom[556] = 0;
     rom[557] = 1;
     rom[558] = 1;
     rom[559] = 1;
     rom[560] = 1;
     rom[561] = 1;
     rom[562] = 1;
     rom[563] = 1;
     rom[564] = 1;
     rom[565] = 1;
     rom[566] = 1;
     rom[567] = 1;
     rom[568] = 0;
     rom[569] = 0;
     rom[570] = 0;
     rom[571] = 0;
     rom[572] = 0;
     rom[573] = 0;
     rom[574] = 0;
     rom[575] = 0;
     rom[576] = 0;
     rom[577] = 0;
     rom[578] = 0;
     rom[579] = 0;
     rom[580] = 0;
     rom[581] = 0;
     rom[582] = 0;
     rom[583] = 1;
     rom[584] = 1;
     rom[585] = 1;
     rom[586] = 1;
     rom[587] = 1;
     rom[588] = 1;
     rom[589] = 1;
     rom[590] = 1;
     rom[591] = 1;
     rom[592] = 1;
     rom[593] = 1;
     rom[594] = 1;
     rom[595] = 1;
     rom[596] = 0;
     rom[597] = 0;
     rom[598] = 0;
     rom[599] = 0;
     rom[600] = 0;
     rom[601] = 0;
     rom[602] = 1;
     rom[603] = 1;
     rom[604] = 1;
     rom[605] = 1;
     rom[606] = 1;
     rom[607] = 1;
     rom[608] = 1;
     rom[609] = 1;
     rom[610] = 1;
     rom[611] = 1;
     rom[612] = 1;
     rom[613] = 1;
     rom[614] = 0;
     rom[615] = 0;
     rom[616] = 0;
     rom[617] = 0;
     rom[618] = 0;
     rom[619] = 0;
     rom[620] = 1;
     rom[621] = 1;
     rom[622] = 1;
     rom[623] = 1;
     rom[624] = 1;
     rom[625] = 1;
     rom[626] = 1;
     rom[627] = 1;
     rom[628] = 1;
     rom[629] = 1;
     rom[630] = 1;
     rom[631] = 1;
     rom[632] = 1;
     rom[633] = 0;
     rom[634] = 0;
     rom[635] = 0;
     rom[636] = 0;
     rom[637] = 0;
     rom[638] = 0;
     rom[639] = 0;
     rom[640] = 0;
     rom[641] = 0;
     rom[642] = 0;
     rom[643] = 0;
     rom[644] = 0;
     rom[645] = 0;
     rom[646] = 0;
     rom[647] = 1;
     rom[648] = 1;
     rom[649] = 1;
     rom[650] = 1;
     rom[651] = 1;
     rom[652] = 1;
     rom[653] = 1;
     rom[654] = 1;
     rom[655] = 1;
     rom[656] = 1;
     rom[657] = 1;
     rom[658] = 1;
     rom[659] = 1;
     rom[660] = 0;
     rom[661] = 0;
     rom[662] = 0;
     rom[663] = 0;
     rom[664] = 0;
     rom[665] = 1;
     rom[666] = 1;
     rom[667] = 1;
     rom[668] = 1;
     rom[669] = 1;
     rom[670] = 1;
     rom[671] = 1;
     rom[672] = 1;
     rom[673] = 1;
     rom[674] = 1;
     rom[675] = 1;
     rom[676] = 1;
     rom[677] = 1;
     rom[678] = 1;
     rom[679] = 0;
     rom[680] = 0;
     rom[681] = 0;
     rom[682] = 0;
     rom[683] = 1;
     rom[684] = 1;
     rom[685] = 1;
     rom[686] = 1;
     rom[687] = 1;
     rom[688] = 1;
     rom[689] = 1;
     rom[690] = 1;
     rom[691] = 1;
     rom[692] = 1;
     rom[693] = 1;
     rom[694] = 1;
     rom[695] = 1;
     rom[696] = 1;
     rom[697] = 0;
     rom[698] = 0;
     rom[699] = 0;
     rom[700] = 0;
     rom[701] = 0;
     rom[702] = 0;
     rom[703] = 0;
     rom[704] = 0;
     rom[705] = 0;
     rom[706] = 0;
     rom[707] = 0;
     rom[708] = 0;
     rom[709] = 0;
     rom[710] = 0;
     rom[711] = 1;
     rom[712] = 1;
     rom[713] = 1;
     rom[714] = 1;
     rom[715] = 1;
     rom[716] = 1;
     rom[717] = 1;
     rom[718] = 1;
     rom[719] = 1;
     rom[720] = 1;
     rom[721] = 1;
     rom[722] = 1;
     rom[723] = 1;
     rom[724] = 1;
     rom[725] = 0;
     rom[726] = 0;
     rom[727] = 0;
     rom[728] = 0;
     rom[729] = 1;
     rom[730] = 1;
     rom[731] = 1;
     rom[732] = 1;
     rom[733] = 1;
     rom[734] = 1;
     rom[735] = 1;
     rom[736] = 1;
     rom[737] = 1;
     rom[738] = 1;
     rom[739] = 1;
     rom[740] = 1;
     rom[741] = 1;
     rom[742] = 1;
     rom[743] = 0;
     rom[744] = 0;
     rom[745] = 0;
     rom[746] = 0;
     rom[747] = 1;
     rom[748] = 1;
     rom[749] = 1;
     rom[750] = 1;
     rom[751] = 1;
     rom[752] = 1;
     rom[753] = 1;
     rom[754] = 1;
     rom[755] = 1;
     rom[756] = 1;
     rom[757] = 1;
     rom[758] = 1;
     rom[759] = 1;
     rom[760] = 1;
     rom[761] = 0;
     rom[762] = 0;
     rom[763] = 0;
     rom[764] = 0;
     rom[765] = 0;
     rom[766] = 0;
     rom[767] = 0;
     rom[768] = 0;
     rom[769] = 0;
     rom[770] = 0;
     rom[771] = 0;
     rom[772] = 0;
     rom[773] = 0;
     rom[774] = 1;
     rom[775] = 1;
     rom[776] = 1;
     rom[777] = 1;
     rom[778] = 1;
     rom[779] = 1;
     rom[780] = 1;
     rom[781] = 1;
     rom[782] = 1;
     rom[783] = 1;
     rom[784] = 1;
     rom[785] = 1;
     rom[786] = 1;
     rom[787] = 1;
     rom[788] = 1;
     rom[789] = 0;
     rom[790] = 0;
     rom[791] = 0;
     rom[792] = 0;
     rom[793] = 1;
     rom[794] = 1;
     rom[795] = 1;
     rom[796] = 1;
     rom[797] = 1;
     rom[798] = 1;
     rom[799] = 1;
     rom[800] = 1;
     rom[801] = 1;
     rom[802] = 1;
     rom[803] = 1;
     rom[804] = 1;
     rom[805] = 1;
     rom[806] = 1;
     rom[807] = 0;
     rom[808] = 0;
     rom[809] = 0;
     rom[810] = 0;
     rom[811] = 1;
     rom[812] = 1;
     rom[813] = 1;
     rom[814] = 1;
     rom[815] = 1;
     rom[816] = 1;
     rom[817] = 1;
     rom[818] = 1;
     rom[819] = 1;
     rom[820] = 1;
     rom[821] = 1;
     rom[822] = 1;
     rom[823] = 1;
     rom[824] = 1;
     rom[825] = 1;
     rom[826] = 0;
     rom[827] = 0;
     rom[828] = 0;
     rom[829] = 0;
     rom[830] = 0;
     rom[831] = 0;
     rom[832] = 0;
     rom[833] = 0;
     rom[834] = 0;
     rom[835] = 0;
     rom[836] = 0;
     rom[837] = 0;
     rom[838] = 1;
     rom[839] = 1;
     rom[840] = 1;
     rom[841] = 1;
     rom[842] = 1;
     rom[843] = 1;
     rom[844] = 1;
     rom[845] = 1;
     rom[846] = 1;
     rom[847] = 1;
     rom[848] = 1;
     rom[849] = 1;
     rom[850] = 1;
     rom[851] = 1;
     rom[852] = 1;
     rom[853] = 0;
     rom[854] = 0;
     rom[855] = 0;
     rom[856] = 0;
     rom[857] = 1;
     rom[858] = 1;
     rom[859] = 1;
     rom[860] = 1;
     rom[861] = 1;
     rom[862] = 1;
     rom[863] = 1;
     rom[864] = 1;
     rom[865] = 1;
     rom[866] = 1;
     rom[867] = 1;
     rom[868] = 1;
     rom[869] = 1;
     rom[870] = 1;
     rom[871] = 0;
     rom[872] = 0;
     rom[873] = 0;
     rom[874] = 0;
     rom[875] = 1;
     rom[876] = 1;
     rom[877] = 1;
     rom[878] = 1;
     rom[879] = 1;
     rom[880] = 1;
     rom[881] = 1;
     rom[882] = 1;
     rom[883] = 1;
     rom[884] = 1;
     rom[885] = 1;
     rom[886] = 1;
     rom[887] = 1;
     rom[888] = 1;
     rom[889] = 1;
     rom[890] = 0;
     rom[891] = 0;
     rom[892] = 0;
     rom[893] = 0;
     rom[894] = 0;
     rom[895] = 0;
     rom[896] = 0;
     rom[897] = 0;
     rom[898] = 0;
     rom[899] = 0;
     rom[900] = 0;
     rom[901] = 0;
     rom[902] = 1;
     rom[903] = 1;
     rom[904] = 1;
     rom[905] = 1;
     rom[906] = 1;
     rom[907] = 1;
     rom[908] = 1;
     rom[909] = 1;
     rom[910] = 1;
     rom[911] = 1;
     rom[912] = 1;
     rom[913] = 1;
     rom[914] = 1;
     rom[915] = 1;
     rom[916] = 1;
     rom[917] = 0;
     rom[918] = 0;
     rom[919] = 0;
     rom[920] = 0;
     rom[921] = 1;
     rom[922] = 1;
     rom[923] = 1;
     rom[924] = 1;
     rom[925] = 1;
     rom[926] = 1;
     rom[927] = 1;
     rom[928] = 1;
     rom[929] = 1;
     rom[930] = 1;
     rom[931] = 1;
     rom[932] = 1;
     rom[933] = 1;
     rom[934] = 1;
     rom[935] = 0;
     rom[936] = 0;
     rom[937] = 0;
     rom[938] = 0;
     rom[939] = 1;
     rom[940] = 1;
     rom[941] = 1;
     rom[942] = 1;
     rom[943] = 1;
     rom[944] = 1;
     rom[945] = 1;
     rom[946] = 1;
     rom[947] = 1;
     rom[948] = 1;
     rom[949] = 1;
     rom[950] = 1;
     rom[951] = 1;
     rom[952] = 1;
     rom[953] = 1;
     rom[954] = 0;
     rom[955] = 0;
     rom[956] = 0;
     rom[957] = 0;
     rom[958] = 0;
     rom[959] = 0;
     rom[960] = 0;
     rom[961] = 0;
     rom[962] = 0;
     rom[963] = 0;
     rom[964] = 0;
     rom[965] = 0;
     rom[966] = 0;
     rom[967] = 1;
     rom[968] = 1;
     rom[969] = 1;
     rom[970] = 1;
     rom[971] = 1;
     rom[972] = 1;
     rom[973] = 1;
     rom[974] = 1;
     rom[975] = 1;
     rom[976] = 1;
     rom[977] = 1;
     rom[978] = 1;
     rom[979] = 1;
     rom[980] = 1;
     rom[981] = 0;
     rom[982] = 0;
     rom[983] = 0;
     rom[984] = 0;
     rom[985] = 1;
     rom[986] = 1;
     rom[987] = 1;
     rom[988] = 1;
     rom[989] = 1;
     rom[990] = 1;
     rom[991] = 1;
     rom[992] = 1;
     rom[993] = 1;
     rom[994] = 1;
     rom[995] = 1;
     rom[996] = 1;
     rom[997] = 1;
     rom[998] = 1;
     rom[999] = 0;
     rom[1000] = 0;
     rom[1001] = 0;
     rom[1002] = 0;
     rom[1003] = 1;
     rom[1004] = 1;
     rom[1005] = 1;
     rom[1006] = 1;
     rom[1007] = 1;
     rom[1008] = 1;
     rom[1009] = 1;
     rom[1010] = 1;
     rom[1011] = 1;
     rom[1012] = 1;
     rom[1013] = 1;
     rom[1014] = 1;
     rom[1015] = 1;
     rom[1016] = 1;
     rom[1017] = 0;
     rom[1018] = 0;
     rom[1019] = 0;
     rom[1020] = 0;
     rom[1021] = 0;
     rom[1022] = 0;
     rom[1023] = 0;
     rom[1024] = 0;
     rom[1025] = 0;
     rom[1026] = 0;
     rom[1027] = 0;
     rom[1028] = 0;
     rom[1029] = 0;
     rom[1030] = 0;
     rom[1031] = 1;
     rom[1032] = 1;
     rom[1033] = 1;
     rom[1034] = 1;
     rom[1035] = 1;
     rom[1036] = 1;
     rom[1037] = 1;
     rom[1038] = 1;
     rom[1039] = 1;
     rom[1040] = 1;
     rom[1041] = 1;
     rom[1042] = 1;
     rom[1043] = 1;
     rom[1044] = 0;
     rom[1045] = 0;
     rom[1046] = 0;
     rom[1047] = 0;
     rom[1048] = 0;
     rom[1049] = 1;
     rom[1050] = 1;
     rom[1051] = 1;
     rom[1052] = 1;
     rom[1053] = 1;
     rom[1054] = 1;
     rom[1055] = 1;
     rom[1056] = 1;
     rom[1057] = 1;
     rom[1058] = 1;
     rom[1059] = 1;
     rom[1060] = 1;
     rom[1061] = 1;
     rom[1062] = 1;
     rom[1063] = 0;
     rom[1064] = 0;
     rom[1065] = 0;
     rom[1066] = 0;
     rom[1067] = 1;
     rom[1068] = 1;
     rom[1069] = 1;
     rom[1070] = 1;
     rom[1071] = 1;
     rom[1072] = 1;
     rom[1073] = 1;
     rom[1074] = 1;
     rom[1075] = 1;
     rom[1076] = 1;
     rom[1077] = 1;
     rom[1078] = 1;
     rom[1079] = 1;
     rom[1080] = 1;
     rom[1081] = 0;
     rom[1082] = 0;
     rom[1083] = 0;
     rom[1084] = 0;
     rom[1085] = 0;
     rom[1086] = 0;
     rom[1087] = 0;
     rom[1088] = 0;
     rom[1089] = 0;
     rom[1090] = 0;
     rom[1091] = 0;
     rom[1092] = 0;
     rom[1093] = 0;
     rom[1094] = 0;
     rom[1095] = 1;
     rom[1096] = 1;
     rom[1097] = 1;
     rom[1098] = 1;
     rom[1099] = 1;
     rom[1100] = 1;
     rom[1101] = 1;
     rom[1102] = 1;
     rom[1103] = 1;
     rom[1104] = 1;
     rom[1105] = 1;
     rom[1106] = 1;
     rom[1107] = 1;
     rom[1108] = 0;
     rom[1109] = 0;
     rom[1110] = 0;
     rom[1111] = 0;
     rom[1112] = 0;
     rom[1113] = 0;
     rom[1114] = 1;
     rom[1115] = 1;
     rom[1116] = 1;
     rom[1117] = 1;
     rom[1118] = 1;
     rom[1119] = 1;
     rom[1120] = 1;
     rom[1121] = 1;
     rom[1122] = 1;
     rom[1123] = 1;
     rom[1124] = 1;
     rom[1125] = 1;
     rom[1126] = 0;
     rom[1127] = 0;
     rom[1128] = 0;
     rom[1129] = 0;
     rom[1130] = 0;
     rom[1131] = 0;
     rom[1132] = 1;
     rom[1133] = 1;
     rom[1134] = 1;
     rom[1135] = 1;
     rom[1136] = 1;
     rom[1137] = 1;
     rom[1138] = 1;
     rom[1139] = 1;
     rom[1140] = 1;
     rom[1141] = 1;
     rom[1142] = 1;
     rom[1143] = 1;
     rom[1144] = 0;
     rom[1145] = 0;
     rom[1146] = 0;
     rom[1147] = 0;
     rom[1148] = 0;
     rom[1149] = 0;
     rom[1150] = 0;
     rom[1151] = 0;
     rom[1152] = 0;
     rom[1153] = 0;
     rom[1154] = 0;
     rom[1155] = 0;
     rom[1156] = 0;
     rom[1157] = 0;
     rom[1158] = 0;
     rom[1159] = 0;
     rom[1160] = 1;
     rom[1161] = 1;
     rom[1162] = 1;
     rom[1163] = 1;
     rom[1164] = 1;
     rom[1165] = 1;
     rom[1166] = 1;
     rom[1167] = 1;
     rom[1168] = 1;
     rom[1169] = 1;
     rom[1170] = 1;
     rom[1171] = 0;
     rom[1172] = 0;
     rom[1173] = 0;
     rom[1174] = 0;
     rom[1175] = 0;
     rom[1176] = 0;
     rom[1177] = 0;
     rom[1178] = 1;
     rom[1179] = 1;
     rom[1180] = 1;
     rom[1181] = 1;
     rom[1182] = 1;
     rom[1183] = 1;
     rom[1184] = 1;
     rom[1185] = 1;
     rom[1186] = 1;
     rom[1187] = 1;
     rom[1188] = 1;
     rom[1189] = 0;
     rom[1190] = 0;
     rom[1191] = 0;
     rom[1192] = 0;
     rom[1193] = 0;
     rom[1194] = 0;
     rom[1195] = 0;
     rom[1196] = 0;
     rom[1197] = 1;
     rom[1198] = 1;
     rom[1199] = 1;
     rom[1200] = 1;
     rom[1201] = 1;
     rom[1202] = 1;
     rom[1203] = 1;
     rom[1204] = 1;
     rom[1205] = 1;
     rom[1206] = 1;
     rom[1207] = 1;
     rom[1208] = 0;
     rom[1209] = 0;
     rom[1210] = 0;
     rom[1211] = 0;
     rom[1212] = 0;
     rom[1213] = 0;
     rom[1214] = 0;
     rom[1215] = 0;
     rom[1216] = 0;
     rom[1217] = 0;
     rom[1218] = 0;
     rom[1219] = 0;
     rom[1220] = 0;
     rom[1221] = 0;
     rom[1222] = 0;
     rom[1223] = 0;
     rom[1224] = 0;
     rom[1225] = 1;
     rom[1226] = 1;
     rom[1227] = 1;
     rom[1228] = 1;
     rom[1229] = 1;
     rom[1230] = 1;
     rom[1231] = 1;
     rom[1232] = 1;
     rom[1233] = 1;
     rom[1234] = 0;
     rom[1235] = 0;
     rom[1236] = 0;
     rom[1237] = 0;
     rom[1238] = 0;
     rom[1239] = 0;
     rom[1240] = 0;
     rom[1241] = 0;
     rom[1242] = 0;
     rom[1243] = 0;
     rom[1244] = 1;
     rom[1245] = 1;
     rom[1246] = 1;
     rom[1247] = 1;
     rom[1248] = 1;
     rom[1249] = 1;
     rom[1250] = 1;
     rom[1251] = 1;
     rom[1252] = 0;
     rom[1253] = 0;
     rom[1254] = 0;
     rom[1255] = 0;
     rom[1256] = 0;
     rom[1257] = 0;
     rom[1258] = 0;
     rom[1259] = 0;
     rom[1260] = 0;
     rom[1261] = 0;
     rom[1262] = 1;
     rom[1263] = 1;
     rom[1264] = 1;
     rom[1265] = 1;
     rom[1266] = 1;
     rom[1267] = 1;
     rom[1268] = 1;
     rom[1269] = 1;
     rom[1270] = 1;
     rom[1271] = 0;
     rom[1272] = 0;
     rom[1273] = 0;
     rom[1274] = 0;
     rom[1275] = 0;
     rom[1276] = 0;
     rom[1277] = 0;
     rom[1278] = 0;
     rom[1279] = 0;
     rom[1280] = 0;
     rom[1281] = 0;
     rom[1282] = 0;
     rom[1283] = 0;
     rom[1284] = 0;
     rom[1285] = 0;
     rom[1286] = 0;
     rom[1287] = 0;
     rom[1288] = 0;
     rom[1289] = 0;
     rom[1290] = 0;
     rom[1291] = 1;
     rom[1292] = 1;
     rom[1293] = 1;
     rom[1294] = 1;
     rom[1295] = 1;
     rom[1296] = 0;
     rom[1297] = 0;
     rom[1298] = 0;
     rom[1299] = 0;
     rom[1300] = 0;
     rom[1301] = 0;
     rom[1302] = 0;
     rom[1303] = 0;
     rom[1304] = 0;
     rom[1305] = 0;
     rom[1306] = 0;
     rom[1307] = 0;
     rom[1308] = 0;
     rom[1309] = 0;
     rom[1310] = 1;
     rom[1311] = 1;
     rom[1312] = 1;
     rom[1313] = 1;
     rom[1314] = 0;
     rom[1315] = 0;
     rom[1316] = 0;
     rom[1317] = 0;
     rom[1318] = 0;
     rom[1319] = 0;
     rom[1320] = 0;
     rom[1321] = 0;
     rom[1322] = 0;
     rom[1323] = 0;
     rom[1324] = 0;
     rom[1325] = 0;
     rom[1326] = 0;
     rom[1327] = 0;
     rom[1328] = 1;
     rom[1329] = 1;
     rom[1330] = 1;
     rom[1331] = 1;
     rom[1332] = 1;
     rom[1333] = 0;
     rom[1334] = 0;
     rom[1335] = 0;
     rom[1336] = 0;
     rom[1337] = 0;
     rom[1338] = 0;
     rom[1339] = 0;
     rom[1340] = 0;
     rom[1341] = 0;
     rom[1342] = 0;
     rom[1343] = 0;
     rom[1344] = 0;
     rom[1345] = 0;
     rom[1346] = 0;
     rom[1347] = 0;
     rom[1348] = 0;
     rom[1349] = 0;
     rom[1350] = 0;
     rom[1351] = 0;
     rom[1352] = 0;
     rom[1353] = 0;
     rom[1354] = 0;
     rom[1355] = 0;
     rom[1356] = 0;
     rom[1357] = 0;
     rom[1358] = 0;
     rom[1359] = 0;
     rom[1360] = 0;
     rom[1361] = 0;
     rom[1362] = 0;
     rom[1363] = 0;
     rom[1364] = 0;
     rom[1365] = 0;
     rom[1366] = 0;
     rom[1367] = 0;
     rom[1368] = 0;
     rom[1369] = 0;
     rom[1370] = 0;
     rom[1371] = 0;
     rom[1372] = 0;
     rom[1373] = 0;
     rom[1374] = 0;
     rom[1375] = 0;
     rom[1376] = 0;
     rom[1377] = 0;
     rom[1378] = 0;
     rom[1379] = 0;
     rom[1380] = 0;
     rom[1381] = 0;
     rom[1382] = 0;
     rom[1383] = 0;
     rom[1384] = 0;
     rom[1385] = 0;
     rom[1386] = 0;
     rom[1387] = 0;
     rom[1388] = 0;
     rom[1389] = 0;
     rom[1390] = 0;
     rom[1391] = 0;
     rom[1392] = 0;
     rom[1393] = 0;
     rom[1394] = 0;
     rom[1395] = 0;
     rom[1396] = 0;
     rom[1397] = 0;
     rom[1398] = 0;
     rom[1399] = 0;
     rom[1400] = 0;
     rom[1401] = 0;
     rom[1402] = 0;
     rom[1403] = 0;
     rom[1404] = 0;
     rom[1405] = 0;
     rom[1406] = 0;
     rom[1407] = 0;
     rom[1408] = 0;
     rom[1409] = 0;
     rom[1410] = 0;
     rom[1411] = 0;
     rom[1412] = 0;
     rom[1413] = 0;
     rom[1414] = 0;
     rom[1415] = 0;
     rom[1416] = 0;
     rom[1417] = 0;
     rom[1418] = 0;
     rom[1419] = 0;
     rom[1420] = 0;
     rom[1421] = 0;
     rom[1422] = 0;
     rom[1423] = 0;
     rom[1424] = 0;
     rom[1425] = 0;
     rom[1426] = 0;
     rom[1427] = 0;
     rom[1428] = 0;
     rom[1429] = 0;
     rom[1430] = 0;
     rom[1431] = 0;
     rom[1432] = 0;
     rom[1433] = 0;
     rom[1434] = 0;
     rom[1435] = 0;
     rom[1436] = 0;
     rom[1437] = 0;
     rom[1438] = 0;
     rom[1439] = 0;
     rom[1440] = 0;
     rom[1441] = 0;
     rom[1442] = 0;
     rom[1443] = 0;
     rom[1444] = 0;
     rom[1445] = 0;
     rom[1446] = 0;
     rom[1447] = 0;
     rom[1448] = 0;
     rom[1449] = 0;
     rom[1450] = 0;
     rom[1451] = 0;
     rom[1452] = 0;
     rom[1453] = 0;
     rom[1454] = 0;
     rom[1455] = 0;
     rom[1456] = 0;
     rom[1457] = 0;
     rom[1458] = 0;
     rom[1459] = 0;
     rom[1460] = 0;
     rom[1461] = 0;
     rom[1462] = 0;
     rom[1463] = 0;
     rom[1464] = 0;
     rom[1465] = 0;
     rom[1466] = 0;
     rom[1467] = 0;
     rom[1468] = 0;
     rom[1469] = 0;
     rom[1470] = 0;
     rom[1471] = 0;
     rom[1472] = 0;
     rom[1473] = 0;
     rom[1474] = 0;
     rom[1475] = 0;
     rom[1476] = 0;
     rom[1477] = 0;
     rom[1478] = 0;
     rom[1479] = 0;
     rom[1480] = 0;
     rom[1481] = 0;
     rom[1482] = 0;
     rom[1483] = 0;
     rom[1484] = 0;
     rom[1485] = 0;
     rom[1486] = 0;
     rom[1487] = 0;
     rom[1488] = 0;
     rom[1489] = 0;
     rom[1490] = 0;
     rom[1491] = 0;
     rom[1492] = 0;
     rom[1493] = 0;
     rom[1494] = 0;
     rom[1495] = 0;
     rom[1496] = 0;
     rom[1497] = 0;
     rom[1498] = 0;
     rom[1499] = 0;
     rom[1500] = 0;
     rom[1501] = 0;
     rom[1502] = 0;
     rom[1503] = 0;
     rom[1504] = 0;
     rom[1505] = 0;
     rom[1506] = 0;
     rom[1507] = 0;
     rom[1508] = 0;
     rom[1509] = 0;
     rom[1510] = 0;
     rom[1511] = 0;
     rom[1512] = 0;
     rom[1513] = 0;
     rom[1514] = 0;
     rom[1515] = 0;
     rom[1516] = 0;
     rom[1517] = 0;
     rom[1518] = 0;
     rom[1519] = 0;
     rom[1520] = 0;
     rom[1521] = 0;
     rom[1522] = 0;
     rom[1523] = 0;
     rom[1524] = 0;
     rom[1525] = 0;
     rom[1526] = 0;
     rom[1527] = 0;
     rom[1528] = 0;
     rom[1529] = 0;
     rom[1530] = 0;
     rom[1531] = 0;
     rom[1532] = 0;
     rom[1533] = 0;
     rom[1534] = 0;
     rom[1535] = 0;
     rom[1536] = 0;
     rom[1537] = 0;
     rom[1538] = 0;
     rom[1539] = 0;
     rom[1540] = 0;
     rom[1541] = 0;
     rom[1542] = 0;
     rom[1543] = 0;
     rom[1544] = 0;
     rom[1545] = 0;
     rom[1546] = 0;
     rom[1547] = 0;
     rom[1548] = 0;
     rom[1549] = 0;
     rom[1550] = 0;
     rom[1551] = 0;
     rom[1552] = 0;
     rom[1553] = 0;
     rom[1554] = 0;
     rom[1555] = 0;
     rom[1556] = 0;
     rom[1557] = 0;
     rom[1558] = 0;
     rom[1559] = 0;
     rom[1560] = 0;
     rom[1561] = 0;
     rom[1562] = 0;
     rom[1563] = 0;
     rom[1564] = 0;
     rom[1565] = 0;
     rom[1566] = 0;
     rom[1567] = 0;
     rom[1568] = 0;
     rom[1569] = 0;
     rom[1570] = 0;
     rom[1571] = 0;
     rom[1572] = 0;
     rom[1573] = 0;
     rom[1574] = 0;
     rom[1575] = 0;
     rom[1576] = 0;
     rom[1577] = 0;
     rom[1578] = 0;
     rom[1579] = 0;
     rom[1580] = 0;
     rom[1581] = 0;
     rom[1582] = 0;
     rom[1583] = 0;
     rom[1584] = 0;
     rom[1585] = 0;
     rom[1586] = 0;
     rom[1587] = 0;
     rom[1588] = 0;
     rom[1589] = 0;
     rom[1590] = 0;
     rom[1591] = 0;
     rom[1592] = 0;
     rom[1593] = 0;
     rom[1594] = 0;
     rom[1595] = 0;
     rom[1596] = 0;
     rom[1597] = 0;
     rom[1598] = 0;
     rom[1599] = 0;
     rom[1600] = 0;
     rom[1601] = 0;
     rom[1602] = 0;
     rom[1603] = 0;
     rom[1604] = 0;
     rom[1605] = 0;
     rom[1606] = 0;
     rom[1607] = 0;
     rom[1608] = 0;
     rom[1609] = 0;
     rom[1610] = 0;
     rom[1611] = 0;
     rom[1612] = 0;
     rom[1613] = 0;
     rom[1614] = 0;
     rom[1615] = 0;
     rom[1616] = 0;
     rom[1617] = 0;
     rom[1618] = 0;
     rom[1619] = 0;
     rom[1620] = 0;
     rom[1621] = 0;
     rom[1622] = 0;
     rom[1623] = 0;
     rom[1624] = 0;
     rom[1625] = 0;
     rom[1626] = 0;
     rom[1627] = 0;
     rom[1628] = 0;
     rom[1629] = 0;
     rom[1630] = 0;
     rom[1631] = 0;
     rom[1632] = 0;
     rom[1633] = 0;
     rom[1634] = 0;
     rom[1635] = 0;
     rom[1636] = 0;
     rom[1637] = 0;
     rom[1638] = 0;
     rom[1639] = 0;
     rom[1640] = 0;
     rom[1641] = 0;
     rom[1642] = 0;
     rom[1643] = 0;
     rom[1644] = 0;
     rom[1645] = 0;
     rom[1646] = 0;
     rom[1647] = 0;
     rom[1648] = 0;
     rom[1649] = 0;
     rom[1650] = 0;
     rom[1651] = 0;
     rom[1652] = 0;
     rom[1653] = 0;
     rom[1654] = 0;
     rom[1655] = 0;
     rom[1656] = 0;
     rom[1657] = 0;
     rom[1658] = 0;
     rom[1659] = 0;
     rom[1660] = 0;
     rom[1661] = 0;
     rom[1662] = 0;
     rom[1663] = 0;
     rom[1664] = 0;
     rom[1665] = 0;
     rom[1666] = 0;
     rom[1667] = 0;
     rom[1668] = 0;
     rom[1669] = 0;
     rom[1670] = 0;
     rom[1671] = 0;
     rom[1672] = 0;
     rom[1673] = 0;
     rom[1674] = 0;
     rom[1675] = 0;
     rom[1676] = 0;
     rom[1677] = 0;
     rom[1678] = 0;
     rom[1679] = 0;
     rom[1680] = 0;
     rom[1681] = 0;
     rom[1682] = 0;
     rom[1683] = 0;
     rom[1684] = 0;
     rom[1685] = 0;
     rom[1686] = 0;
     rom[1687] = 0;
     rom[1688] = 0;
     rom[1689] = 0;
     rom[1690] = 0;
     rom[1691] = 0;
     rom[1692] = 0;
     rom[1693] = 0;
     rom[1694] = 0;
     rom[1695] = 0;
     rom[1696] = 0;
     rom[1697] = 0;
     rom[1698] = 0;
     rom[1699] = 0;
     rom[1700] = 0;
     rom[1701] = 0;
     rom[1702] = 0;
     rom[1703] = 0;
     rom[1704] = 0;
     rom[1705] = 0;
     rom[1706] = 0;
     rom[1707] = 0;
     rom[1708] = 0;
     rom[1709] = 0;
     rom[1710] = 0;
     rom[1711] = 0;
     rom[1712] = 0;
     rom[1713] = 0;
     rom[1714] = 0;
     rom[1715] = 0;
     rom[1716] = 0;
     rom[1717] = 0;
     rom[1718] = 0;
     rom[1719] = 0;
     rom[1720] = 0;
     rom[1721] = 0;
     rom[1722] = 0;
     rom[1723] = 0;
     rom[1724] = 0;
     rom[1725] = 0;
     rom[1726] = 0;
     rom[1727] = 0;
     rom[1728] = 0;
     rom[1729] = 0;
     rom[1730] = 0;
     rom[1731] = 0;
     rom[1732] = 0;
     rom[1733] = 0;
     rom[1734] = 0;
     rom[1735] = 0;
     rom[1736] = 0;
     rom[1737] = 0;
     rom[1738] = 0;
     rom[1739] = 0;
     rom[1740] = 0;
     rom[1741] = 0;
     rom[1742] = 0;
     rom[1743] = 0;
     rom[1744] = 0;
     rom[1745] = 0;
     rom[1746] = 0;
     rom[1747] = 0;
     rom[1748] = 0;
     rom[1749] = 0;
     rom[1750] = 0;
     rom[1751] = 0;
     rom[1752] = 0;
     rom[1753] = 0;
     rom[1754] = 0;
     rom[1755] = 0;
     rom[1756] = 0;
     rom[1757] = 0;
     rom[1758] = 0;
     rom[1759] = 0;
     rom[1760] = 0;
     rom[1761] = 0;
     rom[1762] = 0;
     rom[1763] = 0;
     rom[1764] = 0;
     rom[1765] = 0;
     rom[1766] = 0;
     rom[1767] = 0;
     rom[1768] = 0;
     rom[1769] = 0;
     rom[1770] = 0;
     rom[1771] = 0;
     rom[1772] = 0;
     rom[1773] = 0;
     rom[1774] = 0;
     rom[1775] = 0;
     rom[1776] = 0;
     rom[1777] = 0;
     rom[1778] = 0;
     rom[1779] = 0;
     rom[1780] = 0;
     rom[1781] = 0;
     rom[1782] = 0;
     rom[1783] = 0;
     rom[1784] = 0;
     rom[1785] = 0;
     rom[1786] = 0;
     rom[1787] = 0;
     rom[1788] = 0;
     rom[1789] = 0;
     rom[1790] = 0;
     rom[1791] = 0;
     rom[1792] = 0;
     rom[1793] = 0;
     rom[1794] = 0;
     rom[1795] = 0;
     rom[1796] = 0;
     rom[1797] = 0;
     rom[1798] = 0;
     rom[1799] = 0;
     rom[1800] = 0;
     rom[1801] = 0;
     rom[1802] = 0;
     rom[1803] = 0;
     rom[1804] = 0;
     rom[1805] = 0;
     rom[1806] = 0;
     rom[1807] = 0;
     rom[1808] = 0;
     rom[1809] = 0;
     rom[1810] = 0;
     rom[1811] = 0;
     rom[1812] = 0;
     rom[1813] = 0;
     rom[1814] = 0;
     rom[1815] = 0;
     rom[1816] = 0;
     rom[1817] = 0;
     rom[1818] = 0;
     rom[1819] = 0;
     rom[1820] = 0;
     rom[1821] = 0;
     rom[1822] = 0;
     rom[1823] = 0;
     rom[1824] = 0;
     rom[1825] = 0;
     rom[1826] = 0;
     rom[1827] = 0;
     rom[1828] = 0;
     rom[1829] = 0;
     rom[1830] = 0;
     rom[1831] = 0;
     rom[1832] = 0;
     rom[1833] = 0;
     rom[1834] = 0;
     rom[1835] = 0;
     rom[1836] = 0;
     rom[1837] = 0;
     rom[1838] = 0;
     rom[1839] = 0;
     rom[1840] = 0;
     rom[1841] = 0;
     rom[1842] = 0;
     rom[1843] = 0;
     rom[1844] = 0;
     rom[1845] = 0;
     rom[1846] = 0;
     rom[1847] = 0;
     rom[1848] = 0;
     rom[1849] = 0;
     rom[1850] = 0;
     rom[1851] = 0;
     rom[1852] = 0;
     rom[1853] = 0;
     rom[1854] = 0;
     rom[1855] = 0;
     rom[1856] = 0;
     rom[1857] = 0;
     rom[1858] = 0;
     rom[1859] = 0;
     rom[1860] = 0;
     rom[1861] = 0;
     rom[1862] = 0;
     rom[1863] = 0;
     rom[1864] = 0;
     rom[1865] = 0;
     rom[1866] = 0;
     rom[1867] = 0;
     rom[1868] = 0;
     rom[1869] = 0;
     rom[1870] = 0;
     rom[1871] = 0;
     rom[1872] = 0;
     rom[1873] = 0;
     rom[1874] = 0;
     rom[1875] = 0;
     rom[1876] = 0;
     rom[1877] = 0;
     rom[1878] = 0;
     rom[1879] = 0;
     rom[1880] = 0;
     rom[1881] = 0;
     rom[1882] = 0;
     rom[1883] = 0;
     rom[1884] = 0;
     rom[1885] = 0;
     rom[1886] = 0;
     rom[1887] = 0;
     rom[1888] = 0;
     rom[1889] = 0;
     rom[1890] = 0;
     rom[1891] = 0;
     rom[1892] = 0;
     rom[1893] = 0;
     rom[1894] = 0;
     rom[1895] = 0;
     rom[1896] = 0;
     rom[1897] = 0;
     rom[1898] = 0;
     rom[1899] = 0;
     rom[1900] = 0;
     rom[1901] = 0;
     rom[1902] = 0;
     rom[1903] = 0;
     rom[1904] = 0;
     rom[1905] = 0;
     rom[1906] = 0;
     rom[1907] = 0;
     rom[1908] = 0;
     rom[1909] = 0;
     rom[1910] = 0;
     rom[1911] = 0;
     rom[1912] = 0;
     rom[1913] = 0;
     rom[1914] = 0;
     rom[1915] = 0;
     rom[1916] = 0;
     rom[1917] = 0;
     rom[1918] = 0;
     rom[1919] = 0;
     rom[1920] = 0;
     rom[1921] = 0;
     rom[1922] = 0;
     rom[1923] = 0;
     rom[1924] = 0;
     rom[1925] = 0;
     rom[1926] = 0;
     rom[1927] = 0;
     rom[1928] = 0;
     rom[1929] = 0;
     rom[1930] = 0;
     rom[1931] = 0;
     rom[1932] = 0;
     rom[1933] = 0;
     rom[1934] = 0;
     rom[1935] = 0;
     rom[1936] = 0;
     rom[1937] = 0;
     rom[1938] = 0;
     rom[1939] = 0;
     rom[1940] = 0;
     rom[1941] = 0;
     rom[1942] = 0;
     rom[1943] = 0;
     rom[1944] = 0;
     rom[1945] = 0;
     rom[1946] = 0;
     rom[1947] = 0;
     rom[1948] = 0;
     rom[1949] = 0;
     rom[1950] = 0;
     rom[1951] = 0;
     rom[1952] = 0;
     rom[1953] = 0;
     rom[1954] = 0;
     rom[1955] = 0;
     rom[1956] = 0;
     rom[1957] = 0;
     rom[1958] = 0;
     rom[1959] = 0;
     rom[1960] = 0;
     rom[1961] = 0;
     rom[1962] = 0;
     rom[1963] = 0;
     rom[1964] = 0;
     rom[1965] = 0;
     rom[1966] = 0;
     rom[1967] = 0;
     rom[1968] = 0;
     rom[1969] = 0;
     rom[1970] = 0;
     rom[1971] = 0;
     rom[1972] = 0;
     rom[1973] = 0;
     rom[1974] = 0;
     rom[1975] = 0;
     rom[1976] = 0;
     rom[1977] = 0;
     rom[1978] = 0;
     rom[1979] = 0;
     rom[1980] = 0;
     rom[1981] = 0;
     rom[1982] = 0;
     rom[1983] = 0;
     rom[1984] = 0;
     rom[1985] = 0;
     rom[1986] = 0;
     rom[1987] = 0;
     rom[1988] = 0;
     rom[1989] = 0;
     rom[1990] = 0;
     rom[1991] = 0;
     rom[1992] = 0;
     rom[1993] = 0;
     rom[1994] = 0;
     rom[1995] = 0;
     rom[1996] = 0;
     rom[1997] = 0;
     rom[1998] = 0;
     rom[1999] = 0;
     rom[2000] = 0;
     rom[2001] = 0;
     rom[2002] = 0;
     rom[2003] = 0;
     rom[2004] = 0;
     rom[2005] = 0;
     rom[2006] = 0;
     rom[2007] = 0;
     rom[2008] = 0;
     rom[2009] = 0;
     rom[2010] = 0;
     rom[2011] = 0;
     rom[2012] = 0;
     rom[2013] = 0;
     rom[2014] = 0;
     rom[2015] = 0;
     rom[2016] = 0;
     rom[2017] = 0;
     rom[2018] = 0;
     rom[2019] = 0;
     rom[2020] = 0;
     rom[2021] = 0;
     rom[2022] = 0;
     rom[2023] = 0;
     rom[2024] = 0;
     rom[2025] = 0;
     rom[2026] = 0;
     rom[2027] = 0;
     rom[2028] = 0;
     rom[2029] = 0;
     rom[2030] = 0;
     rom[2031] = 0;
     rom[2032] = 0;
     rom[2033] = 0;
     rom[2034] = 0;
     rom[2035] = 0;
     rom[2036] = 0;
     rom[2037] = 0;
     rom[2038] = 0;
     rom[2039] = 0;
     rom[2040] = 0;
     rom[2041] = 0;
     rom[2042] = 0;
     rom[2043] = 0;
     rom[2044] = 0;
     rom[2045] = 0;
     rom[2046] = 0;
     rom[2047] = 0;
     rom[2048] = 0;
     rom[2049] = 0;
     rom[2050] = 0;
     rom[2051] = 0;
     rom[2052] = 0;
     rom[2053] = 0;
     rom[2054] = 0;
     rom[2055] = 0;
     rom[2056] = 0;
     rom[2057] = 0;
     rom[2058] = 0;
     rom[2059] = 0;
     rom[2060] = 0;
     rom[2061] = 0;
     rom[2062] = 0;
     rom[2063] = 0;
     rom[2064] = 0;
     rom[2065] = 0;
     rom[2066] = 0;
     rom[2067] = 0;
     rom[2068] = 0;
     rom[2069] = 0;
     rom[2070] = 0;
     rom[2071] = 0;
     rom[2072] = 0;
     rom[2073] = 0;
     rom[2074] = 0;
     rom[2075] = 0;
     rom[2076] = 0;
     rom[2077] = 0;
     rom[2078] = 0;
     rom[2079] = 0;
     rom[2080] = 0;
     rom[2081] = 0;
     rom[2082] = 0;
     rom[2083] = 0;
     rom[2084] = 0;
     rom[2085] = 0;
     rom[2086] = 0;
     rom[2087] = 0;
     rom[2088] = 0;
     rom[2089] = 0;
     rom[2090] = 0;
     rom[2091] = 0;
     rom[2092] = 0;
     rom[2093] = 0;
     rom[2094] = 0;
     rom[2095] = 0;
     rom[2096] = 0;
     rom[2097] = 0;
     rom[2098] = 0;
     rom[2099] = 0;
     rom[2100] = 0;
     rom[2101] = 0;
     rom[2102] = 0;
     rom[2103] = 0;
     rom[2104] = 0;
     rom[2105] = 0;
     rom[2106] = 0;
     rom[2107] = 0;
     rom[2108] = 0;
     rom[2109] = 0;
     rom[2110] = 0;
     rom[2111] = 0;
     rom[2112] = 0;
     rom[2113] = 0;
     rom[2114] = 0;
     rom[2115] = 0;
     rom[2116] = 0;
     rom[2117] = 0;
     rom[2118] = 0;
     rom[2119] = 0;
     rom[2120] = 0;
     rom[2121] = 0;
     rom[2122] = 0;
     rom[2123] = 0;
     rom[2124] = 0;
     rom[2125] = 0;
     rom[2126] = 0;
     rom[2127] = 0;
     rom[2128] = 0;
     rom[2129] = 0;
     rom[2130] = 0;
     rom[2131] = 0;
     rom[2132] = 0;
     rom[2133] = 0;
     rom[2134] = 0;
     rom[2135] = 0;
     rom[2136] = 0;
     rom[2137] = 0;
     rom[2138] = 0;
     rom[2139] = 0;
     rom[2140] = 0;
     rom[2141] = 0;
     rom[2142] = 0;
     rom[2143] = 0;
     rom[2144] = 0;
     rom[2145] = 0;
     rom[2146] = 0;
     rom[2147] = 0;
     rom[2148] = 0;
     rom[2149] = 0;
     rom[2150] = 0;
     rom[2151] = 0;
     rom[2152] = 0;
     rom[2153] = 0;
     rom[2154] = 0;
     rom[2155] = 0;
     rom[2156] = 0;
     rom[2157] = 0;
     rom[2158] = 0;
     rom[2159] = 0;
     rom[2160] = 0;
     rom[2161] = 0;
     rom[2162] = 0;
     rom[2163] = 0;
     rom[2164] = 0;
     rom[2165] = 0;
     rom[2166] = 0;
     rom[2167] = 0;
     rom[2168] = 0;
     rom[2169] = 0;
     rom[2170] = 0;
     rom[2171] = 0;
     rom[2172] = 0;
     rom[2173] = 0;
     rom[2174] = 0;
     rom[2175] = 0;
     rom[2176] = 0;
     rom[2177] = 0;
     rom[2178] = 0;
     rom[2179] = 0;
     rom[2180] = 0;
     rom[2181] = 0;
     rom[2182] = 0;
     rom[2183] = 0;
     rom[2184] = 0;
     rom[2185] = 0;
     rom[2186] = 0;
     rom[2187] = 0;
     rom[2188] = 0;
     rom[2189] = 0;
     rom[2190] = 0;
     rom[2191] = 0;
     rom[2192] = 0;
     rom[2193] = 0;
     rom[2194] = 0;
     rom[2195] = 0;
     rom[2196] = 0;
     rom[2197] = 0;
     rom[2198] = 0;
     rom[2199] = 0;
     rom[2200] = 0;
     rom[2201] = 0;
     rom[2202] = 0;
     rom[2203] = 0;
     rom[2204] = 0;
     rom[2205] = 0;
     rom[2206] = 0;
     rom[2207] = 0;
     rom[2208] = 0;
     rom[2209] = 0;
     rom[2210] = 0;
     rom[2211] = 0;
     rom[2212] = 0;
     rom[2213] = 0;
     rom[2214] = 0;
     rom[2215] = 0;
     rom[2216] = 0;
     rom[2217] = 0;
     rom[2218] = 0;
     rom[2219] = 0;
     rom[2220] = 0;
     rom[2221] = 0;
     rom[2222] = 0;
     rom[2223] = 0;
     rom[2224] = 0;
     rom[2225] = 0;
     rom[2226] = 0;
     rom[2227] = 0;
     rom[2228] = 0;
     rom[2229] = 0;
     rom[2230] = 0;
     rom[2231] = 0;
     rom[2232] = 0;
     rom[2233] = 0;
     rom[2234] = 0;
     rom[2235] = 0;
     rom[2236] = 0;
     rom[2237] = 0;
     rom[2238] = 0;
     rom[2239] = 0;
     rom[2240] = 0;
     rom[2241] = 0;
     rom[2242] = 0;
     rom[2243] = 0;
     rom[2244] = 0;
     rom[2245] = 0;
     rom[2246] = 0;
     rom[2247] = 0;
     rom[2248] = 0;
     rom[2249] = 0;
     rom[2250] = 0;
     rom[2251] = 0;
     rom[2252] = 0;
     rom[2253] = 0;
     rom[2254] = 0;
     rom[2255] = 0;
     rom[2256] = 0;
     rom[2257] = 0;
     rom[2258] = 0;
     rom[2259] = 0;
     rom[2260] = 0;
     rom[2261] = 0;
     rom[2262] = 0;
     rom[2263] = 0;
     rom[2264] = 0;
     rom[2265] = 0;
     rom[2266] = 0;
     rom[2267] = 0;
     rom[2268] = 0;
     rom[2269] = 0;
     rom[2270] = 0;
     rom[2271] = 0;
     rom[2272] = 0;
     rom[2273] = 0;
     rom[2274] = 0;
     rom[2275] = 0;
     rom[2276] = 0;
     rom[2277] = 0;
     rom[2278] = 0;
     rom[2279] = 0;
     rom[2280] = 0;
     rom[2281] = 0;
     rom[2282] = 0;
     rom[2283] = 0;
     rom[2284] = 0;
     rom[2285] = 0;
     rom[2286] = 0;
     rom[2287] = 0;
     rom[2288] = 0;
     rom[2289] = 0;
     rom[2290] = 0;
     rom[2291] = 0;
     rom[2292] = 0;
     rom[2293] = 0;
     rom[2294] = 0;
     rom[2295] = 0;
     rom[2296] = 0;
     rom[2297] = 0;
     rom[2298] = 0;
     rom[2299] = 0;
     rom[2300] = 0;
     rom[2301] = 0;
     rom[2302] = 0;
     rom[2303] = 0;
     rom[2304] = 0;
     rom[2305] = 0;
     rom[2306] = 0;
     rom[2307] = 0;
     rom[2308] = 0;
     rom[2309] = 0;
     rom[2310] = 0;
     rom[2311] = 0;
     rom[2312] = 0;
     rom[2313] = 0;
     rom[2314] = 0;
     rom[2315] = 0;
     rom[2316] = 0;
     rom[2317] = 0;
     rom[2318] = 0;
     rom[2319] = 0;
     rom[2320] = 0;
     rom[2321] = 0;
     rom[2322] = 0;
     rom[2323] = 0;
     rom[2324] = 0;
     rom[2325] = 0;
     rom[2326] = 0;
     rom[2327] = 0;
     rom[2328] = 0;
     rom[2329] = 0;
     rom[2330] = 0;
     rom[2331] = 0;
     rom[2332] = 0;
     rom[2333] = 0;
     rom[2334] = 0;
     rom[2335] = 0;
     rom[2336] = 0;
     rom[2337] = 0;
     rom[2338] = 0;
     rom[2339] = 0;
     rom[2340] = 0;
     rom[2341] = 0;
     rom[2342] = 0;
     rom[2343] = 0;
     rom[2344] = 0;
     rom[2345] = 0;
     rom[2346] = 0;
     rom[2347] = 0;
     rom[2348] = 0;
     rom[2349] = 0;
     rom[2350] = 0;
     rom[2351] = 0;
     rom[2352] = 0;
     rom[2353] = 0;
     rom[2354] = 0;
     rom[2355] = 0;
     rom[2356] = 0;
     rom[2357] = 0;
     rom[2358] = 0;
     rom[2359] = 0;
     rom[2360] = 0;
     rom[2361] = 0;
     rom[2362] = 0;
     rom[2363] = 0;
     rom[2364] = 0;
     rom[2365] = 0;
     rom[2366] = 0;
     rom[2367] = 0;
     rom[2368] = 0;
     rom[2369] = 0;
     rom[2370] = 0;
     rom[2371] = 0;
     rom[2372] = 0;
     rom[2373] = 0;
     rom[2374] = 0;
     rom[2375] = 0;
     rom[2376] = 0;
     rom[2377] = 0;
     rom[2378] = 0;
     rom[2379] = 0;
     rom[2380] = 0;
     rom[2381] = 0;
     rom[2382] = 0;
     rom[2383] = 0;
     rom[2384] = 0;
     rom[2385] = 0;
     rom[2386] = 0;
     rom[2387] = 0;
     rom[2388] = 0;
     rom[2389] = 0;
     rom[2390] = 0;
     rom[2391] = 0;
     rom[2392] = 0;
     rom[2393] = 0;
     rom[2394] = 0;
     rom[2395] = 0;
     rom[2396] = 0;
     rom[2397] = 0;
     rom[2398] = 0;
     rom[2399] = 0;
     rom[2400] = 0;
     rom[2401] = 0;
     rom[2402] = 0;
     rom[2403] = 0;
     rom[2404] = 0;
     rom[2405] = 0;
     rom[2406] = 0;
     rom[2407] = 0;
     rom[2408] = 0;
     rom[2409] = 0;
     rom[2410] = 0;
     rom[2411] = 0;
     rom[2412] = 0;
     rom[2413] = 0;
     rom[2414] = 0;
     rom[2415] = 0;
     rom[2416] = 0;
     rom[2417] = 0;
     rom[2418] = 0;
     rom[2419] = 0;
     rom[2420] = 0;
     rom[2421] = 0;
     rom[2422] = 0;
     rom[2423] = 0;
     rom[2424] = 0;
     rom[2425] = 0;
     rom[2426] = 0;
     rom[2427] = 0;
     rom[2428] = 0;
     rom[2429] = 0;
     rom[2430] = 0;
     rom[2431] = 0;
     rom[2432] = 0;
     rom[2433] = 0;
     rom[2434] = 0;
     rom[2435] = 0;
     rom[2436] = 0;
     rom[2437] = 0;
     rom[2438] = 0;
     rom[2439] = 0;
     rom[2440] = 0;
     rom[2441] = 0;
     rom[2442] = 0;
     rom[2443] = 0;
     rom[2444] = 0;
     rom[2445] = 0;
     rom[2446] = 0;
     rom[2447] = 0;
     rom[2448] = 0;
     rom[2449] = 0;
     rom[2450] = 0;
     rom[2451] = 0;
     rom[2452] = 0;
     rom[2453] = 0;
     rom[2454] = 0;
     rom[2455] = 0;
     rom[2456] = 0;
     rom[2457] = 0;
     rom[2458] = 0;
     rom[2459] = 0;
     rom[2460] = 0;
     rom[2461] = 0;
     rom[2462] = 0;
     rom[2463] = 0;
     rom[2464] = 0;
     rom[2465] = 0;
     rom[2466] = 0;
     rom[2467] = 0;
     rom[2468] = 0;
     rom[2469] = 0;
     rom[2470] = 0;
     rom[2471] = 0;
     rom[2472] = 0;
     rom[2473] = 0;
     rom[2474] = 0;
     rom[2475] = 0;
     rom[2476] = 0;
     rom[2477] = 0;
     rom[2478] = 0;
     rom[2479] = 0;
     rom[2480] = 0;
     rom[2481] = 0;
     rom[2482] = 0;
     rom[2483] = 0;
     rom[2484] = 0;
     rom[2485] = 0;
     rom[2486] = 0;
     rom[2487] = 0;
     rom[2488] = 0;
     rom[2489] = 0;
     rom[2490] = 0;
     rom[2491] = 0;
     rom[2492] = 0;
     rom[2493] = 0;
     rom[2494] = 0;
     rom[2495] = 0;
     rom[2496] = 0;
     rom[2497] = 0;
     rom[2498] = 0;
     rom[2499] = 0;
     rom[2500] = 0;
     rom[2501] = 0;
     rom[2502] = 0;
     rom[2503] = 0;
     rom[2504] = 0;
     rom[2505] = 0;
     rom[2506] = 0;
     rom[2507] = 0;
     rom[2508] = 0;
     rom[2509] = 0;
     rom[2510] = 0;
     rom[2511] = 0;
     rom[2512] = 0;
     rom[2513] = 0;
     rom[2514] = 0;
     rom[2515] = 0;
     rom[2516] = 0;
     rom[2517] = 0;
     rom[2518] = 0;
     rom[2519] = 0;
     rom[2520] = 0;
     rom[2521] = 0;
     rom[2522] = 0;
     rom[2523] = 0;
     rom[2524] = 0;
     rom[2525] = 0;
     rom[2526] = 0;
     rom[2527] = 0;
     rom[2528] = 0;
     rom[2529] = 0;
     rom[2530] = 0;
     rom[2531] = 0;
     rom[2532] = 0;
     rom[2533] = 0;
     rom[2534] = 0;
     rom[2535] = 0;
     rom[2536] = 0;
     rom[2537] = 0;
     rom[2538] = 0;
     rom[2539] = 0;
     rom[2540] = 0;
     rom[2541] = 0;
     rom[2542] = 0;
     rom[2543] = 0;
     rom[2544] = 0;
     rom[2545] = 0;
     rom[2546] = 0;
     rom[2547] = 0;
     rom[2548] = 0;
     rom[2549] = 0;
     rom[2550] = 0;
     rom[2551] = 0;
     rom[2552] = 0;
     rom[2553] = 0;
     rom[2554] = 0;
     rom[2555] = 0;
     rom[2556] = 0;
     rom[2557] = 0;
     rom[2558] = 0;
     rom[2559] = 0;
     rom[2560] = 0;
     rom[2561] = 0;
     rom[2562] = 0;
     rom[2563] = 0;
     rom[2564] = 0;
     rom[2565] = 0;
     rom[2566] = 0;
     rom[2567] = 0;
     rom[2568] = 0;
     rom[2569] = 0;
     rom[2570] = 0;
     rom[2571] = 0;
     rom[2572] = 0;
     rom[2573] = 0;
     rom[2574] = 0;
     rom[2575] = 0;
     rom[2576] = 0;
     rom[2577] = 0;
     rom[2578] = 0;
     rom[2579] = 0;
     rom[2580] = 0;
     rom[2581] = 0;
     rom[2582] = 0;
     rom[2583] = 0;
     rom[2584] = 0;
     rom[2585] = 0;
     rom[2586] = 0;
     rom[2587] = 0;
     rom[2588] = 0;
     rom[2589] = 0;
     rom[2590] = 0;
     rom[2591] = 0;
     rom[2592] = 0;
     rom[2593] = 0;
     rom[2594] = 0;
     rom[2595] = 0;
     rom[2596] = 0;
     rom[2597] = 0;
     rom[2598] = 0;
     rom[2599] = 0;
     rom[2600] = 0;
     rom[2601] = 0;
     rom[2602] = 0;
     rom[2603] = 0;
     rom[2604] = 0;
     rom[2605] = 0;
     rom[2606] = 0;
     rom[2607] = 0;
     rom[2608] = 0;
     rom[2609] = 0;
     rom[2610] = 0;
     rom[2611] = 0;
     rom[2612] = 0;
     rom[2613] = 0;
     rom[2614] = 0;
     rom[2615] = 0;
     rom[2616] = 0;
     rom[2617] = 0;
     rom[2618] = 0;
     rom[2619] = 0;
     rom[2620] = 0;
     rom[2621] = 0;
     rom[2622] = 0;
     rom[2623] = 0;
     rom[2624] = 0;
     rom[2625] = 0;
     rom[2626] = 0;
     rom[2627] = 0;
     rom[2628] = 0;
     rom[2629] = 0;
     rom[2630] = 0;
     rom[2631] = 0;
     rom[2632] = 0;
     rom[2633] = 0;
     rom[2634] = 0;
     rom[2635] = 0;
     rom[2636] = 0;
     rom[2637] = 0;
     rom[2638] = 0;
     rom[2639] = 0;
     rom[2640] = 0;
     rom[2641] = 0;
     rom[2642] = 0;
     rom[2643] = 0;
     rom[2644] = 0;
     rom[2645] = 0;
     rom[2646] = 0;
     rom[2647] = 0;
     rom[2648] = 0;
     rom[2649] = 0;
     rom[2650] = 0;
     rom[2651] = 0;
     rom[2652] = 0;
     rom[2653] = 0;
     rom[2654] = 0;
     rom[2655] = 0;
     rom[2656] = 0;
     rom[2657] = 0;
     rom[2658] = 0;
     rom[2659] = 0;
     rom[2660] = 0;
     rom[2661] = 0;
     rom[2662] = 0;
     rom[2663] = 0;
     rom[2664] = 0;
     rom[2665] = 0;
     rom[2666] = 0;
     rom[2667] = 0;
     rom[2668] = 0;
     rom[2669] = 0;
     rom[2670] = 0;
     rom[2671] = 0;
     rom[2672] = 0;
     rom[2673] = 0;
     rom[2674] = 0;
     rom[2675] = 0;
     rom[2676] = 0;
     rom[2677] = 0;
     rom[2678] = 0;
     rom[2679] = 0;
     rom[2680] = 0;
     rom[2681] = 0;
     rom[2682] = 0;
     rom[2683] = 0;
     rom[2684] = 0;
     rom[2685] = 0;
     rom[2686] = 0;
     rom[2687] = 0;
     rom[2688] = 0;
     rom[2689] = 0;
     rom[2690] = 0;
     rom[2691] = 0;
     rom[2692] = 0;
     rom[2693] = 0;
     rom[2694] = 0;
     rom[2695] = 0;
     rom[2696] = 0;
     rom[2697] = 0;
     rom[2698] = 0;
     rom[2699] = 0;
     rom[2700] = 0;
     rom[2701] = 0;
     rom[2702] = 0;
     rom[2703] = 0;
     rom[2704] = 0;
     rom[2705] = 0;
     rom[2706] = 0;
     rom[2707] = 0;
     rom[2708] = 0;
     rom[2709] = 0;
     rom[2710] = 0;
     rom[2711] = 0;
     rom[2712] = 0;
     rom[2713] = 0;
     rom[2714] = 0;
     rom[2715] = 0;
     rom[2716] = 0;
     rom[2717] = 0;
     rom[2718] = 0;
     rom[2719] = 0;
     rom[2720] = 0;
     rom[2721] = 0;
     rom[2722] = 0;
     rom[2723] = 0;
     rom[2724] = 0;
     rom[2725] = 0;
     rom[2726] = 0;
     rom[2727] = 0;
     rom[2728] = 0;
     rom[2729] = 0;
     rom[2730] = 0;
     rom[2731] = 0;
     rom[2732] = 0;
     rom[2733] = 0;
     rom[2734] = 0;
     rom[2735] = 0;
     rom[2736] = 0;
     rom[2737] = 0;
     rom[2738] = 0;
     rom[2739] = 0;
     rom[2740] = 0;
     rom[2741] = 0;
     rom[2742] = 0;
     rom[2743] = 0;
     rom[2744] = 0;
     rom[2745] = 0;
     rom[2746] = 0;
     rom[2747] = 0;
     rom[2748] = 0;
     rom[2749] = 0;
     rom[2750] = 0;
     rom[2751] = 0;
     rom[2752] = 0;
     rom[2753] = 0;
     rom[2754] = 0;
     rom[2755] = 0;
     rom[2756] = 0;
     rom[2757] = 0;
     rom[2758] = 0;
     rom[2759] = 0;
     rom[2760] = 0;
     rom[2761] = 0;
     rom[2762] = 0;
     rom[2763] = 1;
     rom[2764] = 1;
     rom[2765] = 1;
     rom[2766] = 1;
     rom[2767] = 1;
     rom[2768] = 0;
     rom[2769] = 0;
     rom[2770] = 0;
     rom[2771] = 0;
     rom[2772] = 0;
     rom[2773] = 0;
     rom[2774] = 0;
     rom[2775] = 0;
     rom[2776] = 0;
     rom[2777] = 0;
     rom[2778] = 0;
     rom[2779] = 0;
     rom[2780] = 0;
     rom[2781] = 0;
     rom[2782] = 1;
     rom[2783] = 1;
     rom[2784] = 1;
     rom[2785] = 1;
     rom[2786] = 0;
     rom[2787] = 0;
     rom[2788] = 0;
     rom[2789] = 0;
     rom[2790] = 0;
     rom[2791] = 0;
     rom[2792] = 0;
     rom[2793] = 0;
     rom[2794] = 0;
     rom[2795] = 0;
     rom[2796] = 0;
     rom[2797] = 0;
     rom[2798] = 0;
     rom[2799] = 0;
     rom[2800] = 1;
     rom[2801] = 1;
     rom[2802] = 1;
     rom[2803] = 1;
     rom[2804] = 1;
     rom[2805] = 0;
     rom[2806] = 0;
     rom[2807] = 0;
     rom[2808] = 0;
     rom[2809] = 0;
     rom[2810] = 0;
     rom[2811] = 0;
     rom[2812] = 0;
     rom[2813] = 0;
     rom[2814] = 0;
     rom[2815] = 0;
     rom[2816] = 0;
     rom[2817] = 0;
     rom[2818] = 0;
     rom[2819] = 0;
     rom[2820] = 0;
     rom[2821] = 0;
     rom[2822] = 0;
     rom[2823] = 0;
     rom[2824] = 0;
     rom[2825] = 1;
     rom[2826] = 1;
     rom[2827] = 1;
     rom[2828] = 1;
     rom[2829] = 1;
     rom[2830] = 1;
     rom[2831] = 1;
     rom[2832] = 1;
     rom[2833] = 1;
     rom[2834] = 0;
     rom[2835] = 0;
     rom[2836] = 0;
     rom[2837] = 0;
     rom[2838] = 0;
     rom[2839] = 0;
     rom[2840] = 0;
     rom[2841] = 0;
     rom[2842] = 0;
     rom[2843] = 0;
     rom[2844] = 1;
     rom[2845] = 1;
     rom[2846] = 1;
     rom[2847] = 1;
     rom[2848] = 1;
     rom[2849] = 1;
     rom[2850] = 1;
     rom[2851] = 1;
     rom[2852] = 0;
     rom[2853] = 0;
     rom[2854] = 0;
     rom[2855] = 0;
     rom[2856] = 0;
     rom[2857] = 0;
     rom[2858] = 0;
     rom[2859] = 0;
     rom[2860] = 0;
     rom[2861] = 0;
     rom[2862] = 1;
     rom[2863] = 1;
     rom[2864] = 1;
     rom[2865] = 1;
     rom[2866] = 1;
     rom[2867] = 1;
     rom[2868] = 1;
     rom[2869] = 1;
     rom[2870] = 1;
     rom[2871] = 0;
     rom[2872] = 0;
     rom[2873] = 0;
     rom[2874] = 0;
     rom[2875] = 0;
     rom[2876] = 0;
     rom[2877] = 0;
     rom[2878] = 0;
     rom[2879] = 0;
     rom[2880] = 0;
     rom[2881] = 0;
     rom[2882] = 0;
     rom[2883] = 0;
     rom[2884] = 0;
     rom[2885] = 0;
     rom[2886] = 0;
     rom[2887] = 0;
     rom[2888] = 1;
     rom[2889] = 1;
     rom[2890] = 1;
     rom[2891] = 1;
     rom[2892] = 1;
     rom[2893] = 1;
     rom[2894] = 1;
     rom[2895] = 1;
     rom[2896] = 1;
     rom[2897] = 1;
     rom[2898] = 1;
     rom[2899] = 0;
     rom[2900] = 0;
     rom[2901] = 0;
     rom[2902] = 0;
     rom[2903] = 0;
     rom[2904] = 0;
     rom[2905] = 0;
     rom[2906] = 1;
     rom[2907] = 1;
     rom[2908] = 1;
     rom[2909] = 1;
     rom[2910] = 1;
     rom[2911] = 1;
     rom[2912] = 1;
     rom[2913] = 1;
     rom[2914] = 1;
     rom[2915] = 1;
     rom[2916] = 1;
     rom[2917] = 0;
     rom[2918] = 0;
     rom[2919] = 0;
     rom[2920] = 0;
     rom[2921] = 0;
     rom[2922] = 0;
     rom[2923] = 0;
     rom[2924] = 0;
     rom[2925] = 1;
     rom[2926] = 1;
     rom[2927] = 1;
     rom[2928] = 1;
     rom[2929] = 1;
     rom[2930] = 1;
     rom[2931] = 1;
     rom[2932] = 1;
     rom[2933] = 1;
     rom[2934] = 1;
     rom[2935] = 1;
     rom[2936] = 0;
     rom[2937] = 0;
     rom[2938] = 0;
     rom[2939] = 0;
     rom[2940] = 0;
     rom[2941] = 0;
     rom[2942] = 0;
     rom[2943] = 0;
     rom[2944] = 0;
     rom[2945] = 0;
     rom[2946] = 0;
     rom[2947] = 0;
     rom[2948] = 0;
     rom[2949] = 0;
     rom[2950] = 0;
     rom[2951] = 1;
     rom[2952] = 1;
     rom[2953] = 1;
     rom[2954] = 1;
     rom[2955] = 1;
     rom[2956] = 1;
     rom[2957] = 1;
     rom[2958] = 1;
     rom[2959] = 1;
     rom[2960] = 1;
     rom[2961] = 1;
     rom[2962] = 1;
     rom[2963] = 1;
     rom[2964] = 0;
     rom[2965] = 0;
     rom[2966] = 0;
     rom[2967] = 0;
     rom[2968] = 0;
     rom[2969] = 0;
     rom[2970] = 1;
     rom[2971] = 1;
     rom[2972] = 1;
     rom[2973] = 1;
     rom[2974] = 1;
     rom[2975] = 1;
     rom[2976] = 1;
     rom[2977] = 1;
     rom[2978] = 1;
     rom[2979] = 1;
     rom[2980] = 1;
     rom[2981] = 1;
     rom[2982] = 0;
     rom[2983] = 0;
     rom[2984] = 0;
     rom[2985] = 0;
     rom[2986] = 0;
     rom[2987] = 0;
     rom[2988] = 1;
     rom[2989] = 1;
     rom[2990] = 1;
     rom[2991] = 1;
     rom[2992] = 1;
     rom[2993] = 1;
     rom[2994] = 1;
     rom[2995] = 1;
     rom[2996] = 1;
     rom[2997] = 1;
     rom[2998] = 1;
     rom[2999] = 1;
     rom[3000] = 0;
     rom[3001] = 0;
     rom[3002] = 0;
     rom[3003] = 0;
     rom[3004] = 0;
     rom[3005] = 0;
     rom[3006] = 0;
     rom[3007] = 0;
     rom[3008] = 0;
     rom[3009] = 0;
     rom[3010] = 0;
     rom[3011] = 0;
     rom[3012] = 0;
     rom[3013] = 0;
     rom[3014] = 0;
     rom[3015] = 1;
     rom[3016] = 1;
     rom[3017] = 1;
     rom[3018] = 1;
     rom[3019] = 1;
     rom[3020] = 1;
     rom[3021] = 1;
     rom[3022] = 1;
     rom[3023] = 1;
     rom[3024] = 1;
     rom[3025] = 1;
     rom[3026] = 1;
     rom[3027] = 1;
     rom[3028] = 0;
     rom[3029] = 0;
     rom[3030] = 0;
     rom[3031] = 0;
     rom[3032] = 0;
     rom[3033] = 1;
     rom[3034] = 1;
     rom[3035] = 1;
     rom[3036] = 1;
     rom[3037] = 1;
     rom[3038] = 1;
     rom[3039] = 1;
     rom[3040] = 1;
     rom[3041] = 1;
     rom[3042] = 1;
     rom[3043] = 1;
     rom[3044] = 1;
     rom[3045] = 1;
     rom[3046] = 1;
     rom[3047] = 0;
     rom[3048] = 0;
     rom[3049] = 0;
     rom[3050] = 0;
     rom[3051] = 1;
     rom[3052] = 1;
     rom[3053] = 1;
     rom[3054] = 1;
     rom[3055] = 1;
     rom[3056] = 1;
     rom[3057] = 1;
     rom[3058] = 1;
     rom[3059] = 1;
     rom[3060] = 1;
     rom[3061] = 1;
     rom[3062] = 1;
     rom[3063] = 1;
     rom[3064] = 1;
     rom[3065] = 0;
     rom[3066] = 0;
     rom[3067] = 0;
     rom[3068] = 0;
     rom[3069] = 0;
     rom[3070] = 0;
     rom[3071] = 0;
     rom[3072] = 0;
     rom[3073] = 0;
     rom[3074] = 0;
     rom[3075] = 0;
     rom[3076] = 0;
     rom[3077] = 0;
     rom[3078] = 0;
     rom[3079] = 1;
     rom[3080] = 1;
     rom[3081] = 1;
     rom[3082] = 1;
     rom[3083] = 1;
     rom[3084] = 1;
     rom[3085] = 1;
     rom[3086] = 1;
     rom[3087] = 1;
     rom[3088] = 1;
     rom[3089] = 1;
     rom[3090] = 1;
     rom[3091] = 1;
     rom[3092] = 1;
     rom[3093] = 0;
     rom[3094] = 0;
     rom[3095] = 0;
     rom[3096] = 0;
     rom[3097] = 1;
     rom[3098] = 1;
     rom[3099] = 1;
     rom[3100] = 1;
     rom[3101] = 1;
     rom[3102] = 1;
     rom[3103] = 1;
     rom[3104] = 1;
     rom[3105] = 1;
     rom[3106] = 1;
     rom[3107] = 1;
     rom[3108] = 1;
     rom[3109] = 1;
     rom[3110] = 1;
     rom[3111] = 0;
     rom[3112] = 0;
     rom[3113] = 0;
     rom[3114] = 0;
     rom[3115] = 1;
     rom[3116] = 1;
     rom[3117] = 1;
     rom[3118] = 1;
     rom[3119] = 1;
     rom[3120] = 1;
     rom[3121] = 1;
     rom[3122] = 1;
     rom[3123] = 1;
     rom[3124] = 1;
     rom[3125] = 1;
     rom[3126] = 1;
     rom[3127] = 1;
     rom[3128] = 1;
     rom[3129] = 0;
     rom[3130] = 0;
     rom[3131] = 0;
     rom[3132] = 0;
     rom[3133] = 0;
     rom[3134] = 0;
     rom[3135] = 0;
     rom[3136] = 0;
     rom[3137] = 0;
     rom[3138] = 0;
     rom[3139] = 0;
     rom[3140] = 0;
     rom[3141] = 0;
     rom[3142] = 1;
     rom[3143] = 1;
     rom[3144] = 1;
     rom[3145] = 1;
     rom[3146] = 1;
     rom[3147] = 1;
     rom[3148] = 1;
     rom[3149] = 1;
     rom[3150] = 1;
     rom[3151] = 1;
     rom[3152] = 1;
     rom[3153] = 1;
     rom[3154] = 1;
     rom[3155] = 1;
     rom[3156] = 1;
     rom[3157] = 0;
     rom[3158] = 0;
     rom[3159] = 0;
     rom[3160] = 0;
     rom[3161] = 1;
     rom[3162] = 1;
     rom[3163] = 1;
     rom[3164] = 1;
     rom[3165] = 1;
     rom[3166] = 1;
     rom[3167] = 1;
     rom[3168] = 1;
     rom[3169] = 1;
     rom[3170] = 1;
     rom[3171] = 1;
     rom[3172] = 1;
     rom[3173] = 1;
     rom[3174] = 1;
     rom[3175] = 0;
     rom[3176] = 0;
     rom[3177] = 0;
     rom[3178] = 0;
     rom[3179] = 1;
     rom[3180] = 1;
     rom[3181] = 1;
     rom[3182] = 1;
     rom[3183] = 1;
     rom[3184] = 1;
     rom[3185] = 1;
     rom[3186] = 1;
     rom[3187] = 1;
     rom[3188] = 1;
     rom[3189] = 1;
     rom[3190] = 1;
     rom[3191] = 1;
     rom[3192] = 1;
     rom[3193] = 1;
     rom[3194] = 0;
     rom[3195] = 0;
     rom[3196] = 0;
     rom[3197] = 0;
     rom[3198] = 0;
     rom[3199] = 0;
     rom[3200] = 0;
     rom[3201] = 0;
     rom[3202] = 0;
     rom[3203] = 0;
     rom[3204] = 0;
     rom[3205] = 0;
     rom[3206] = 1;
     rom[3207] = 1;
     rom[3208] = 1;
     rom[3209] = 1;
     rom[3210] = 1;
     rom[3211] = 1;
     rom[3212] = 1;
     rom[3213] = 1;
     rom[3214] = 1;
     rom[3215] = 1;
     rom[3216] = 1;
     rom[3217] = 1;
     rom[3218] = 1;
     rom[3219] = 1;
     rom[3220] = 1;
     rom[3221] = 0;
     rom[3222] = 0;
     rom[3223] = 0;
     rom[3224] = 0;
     rom[3225] = 1;
     rom[3226] = 1;
     rom[3227] = 1;
     rom[3228] = 1;
     rom[3229] = 1;
     rom[3230] = 1;
     rom[3231] = 1;
     rom[3232] = 1;
     rom[3233] = 1;
     rom[3234] = 1;
     rom[3235] = 1;
     rom[3236] = 1;
     rom[3237] = 1;
     rom[3238] = 1;
     rom[3239] = 0;
     rom[3240] = 0;
     rom[3241] = 0;
     rom[3242] = 0;
     rom[3243] = 1;
     rom[3244] = 1;
     rom[3245] = 1;
     rom[3246] = 1;
     rom[3247] = 1;
     rom[3248] = 1;
     rom[3249] = 1;
     rom[3250] = 1;
     rom[3251] = 1;
     rom[3252] = 1;
     rom[3253] = 1;
     rom[3254] = 1;
     rom[3255] = 1;
     rom[3256] = 1;
     rom[3257] = 1;
     rom[3258] = 0;
     rom[3259] = 0;
     rom[3260] = 0;
     rom[3261] = 0;
     rom[3262] = 0;
     rom[3263] = 0;
     rom[3264] = 0;
     rom[3265] = 0;
     rom[3266] = 0;
     rom[3267] = 0;
     rom[3268] = 0;
     rom[3269] = 0;
     rom[3270] = 1;
     rom[3271] = 1;
     rom[3272] = 1;
     rom[3273] = 1;
     rom[3274] = 1;
     rom[3275] = 1;
     rom[3276] = 1;
     rom[3277] = 1;
     rom[3278] = 1;
     rom[3279] = 1;
     rom[3280] = 1;
     rom[3281] = 1;
     rom[3282] = 1;
     rom[3283] = 1;
     rom[3284] = 1;
     rom[3285] = 0;
     rom[3286] = 0;
     rom[3287] = 0;
     rom[3288] = 0;
     rom[3289] = 1;
     rom[3290] = 1;
     rom[3291] = 1;
     rom[3292] = 1;
     rom[3293] = 1;
     rom[3294] = 1;
     rom[3295] = 1;
     rom[3296] = 1;
     rom[3297] = 1;
     rom[3298] = 1;
     rom[3299] = 1;
     rom[3300] = 1;
     rom[3301] = 1;
     rom[3302] = 1;
     rom[3303] = 0;
     rom[3304] = 0;
     rom[3305] = 0;
     rom[3306] = 0;
     rom[3307] = 1;
     rom[3308] = 1;
     rom[3309] = 1;
     rom[3310] = 1;
     rom[3311] = 1;
     rom[3312] = 1;
     rom[3313] = 1;
     rom[3314] = 1;
     rom[3315] = 1;
     rom[3316] = 1;
     rom[3317] = 1;
     rom[3318] = 1;
     rom[3319] = 1;
     rom[3320] = 1;
     rom[3321] = 1;
     rom[3322] = 0;
     rom[3323] = 0;
     rom[3324] = 0;
     rom[3325] = 0;
     rom[3326] = 0;
     rom[3327] = 0;
     rom[3328] = 0;
     rom[3329] = 0;
     rom[3330] = 0;
     rom[3331] = 0;
     rom[3332] = 0;
     rom[3333] = 0;
     rom[3334] = 0;
     rom[3335] = 1;
     rom[3336] = 1;
     rom[3337] = 1;
     rom[3338] = 1;
     rom[3339] = 1;
     rom[3340] = 1;
     rom[3341] = 1;
     rom[3342] = 1;
     rom[3343] = 1;
     rom[3344] = 1;
     rom[3345] = 1;
     rom[3346] = 1;
     rom[3347] = 1;
     rom[3348] = 1;
     rom[3349] = 0;
     rom[3350] = 0;
     rom[3351] = 0;
     rom[3352] = 0;
     rom[3353] = 1;
     rom[3354] = 1;
     rom[3355] = 1;
     rom[3356] = 1;
     rom[3357] = 1;
     rom[3358] = 1;
     rom[3359] = 1;
     rom[3360] = 1;
     rom[3361] = 1;
     rom[3362] = 1;
     rom[3363] = 1;
     rom[3364] = 1;
     rom[3365] = 1;
     rom[3366] = 1;
     rom[3367] = 0;
     rom[3368] = 0;
     rom[3369] = 0;
     rom[3370] = 0;
     rom[3371] = 1;
     rom[3372] = 1;
     rom[3373] = 1;
     rom[3374] = 1;
     rom[3375] = 1;
     rom[3376] = 1;
     rom[3377] = 1;
     rom[3378] = 1;
     rom[3379] = 1;
     rom[3380] = 1;
     rom[3381] = 1;
     rom[3382] = 1;
     rom[3383] = 1;
     rom[3384] = 1;
     rom[3385] = 0;
     rom[3386] = 0;
     rom[3387] = 0;
     rom[3388] = 0;
     rom[3389] = 0;
     rom[3390] = 0;
     rom[3391] = 0;
     rom[3392] = 0;
     rom[3393] = 0;
     rom[3394] = 0;
     rom[3395] = 0;
     rom[3396] = 0;
     rom[3397] = 0;
     rom[3398] = 0;
     rom[3399] = 1;
     rom[3400] = 1;
     rom[3401] = 1;
     rom[3402] = 1;
     rom[3403] = 1;
     rom[3404] = 1;
     rom[3405] = 1;
     rom[3406] = 1;
     rom[3407] = 1;
     rom[3408] = 1;
     rom[3409] = 1;
     rom[3410] = 1;
     rom[3411] = 1;
     rom[3412] = 0;
     rom[3413] = 0;
     rom[3414] = 0;
     rom[3415] = 0;
     rom[3416] = 0;
     rom[3417] = 1;
     rom[3418] = 1;
     rom[3419] = 1;
     rom[3420] = 1;
     rom[3421] = 1;
     rom[3422] = 1;
     rom[3423] = 1;
     rom[3424] = 1;
     rom[3425] = 1;
     rom[3426] = 1;
     rom[3427] = 1;
     rom[3428] = 1;
     rom[3429] = 1;
     rom[3430] = 1;
     rom[3431] = 0;
     rom[3432] = 0;
     rom[3433] = 0;
     rom[3434] = 0;
     rom[3435] = 1;
     rom[3436] = 1;
     rom[3437] = 1;
     rom[3438] = 1;
     rom[3439] = 1;
     rom[3440] = 1;
     rom[3441] = 1;
     rom[3442] = 1;
     rom[3443] = 1;
     rom[3444] = 1;
     rom[3445] = 1;
     rom[3446] = 1;
     rom[3447] = 1;
     rom[3448] = 1;
     rom[3449] = 0;
     rom[3450] = 0;
     rom[3451] = 0;
     rom[3452] = 0;
     rom[3453] = 0;
     rom[3454] = 0;
     rom[3455] = 0;
     rom[3456] = 0;
     rom[3457] = 0;
     rom[3458] = 0;
     rom[3459] = 0;
     rom[3460] = 0;
     rom[3461] = 0;
     rom[3462] = 0;
     rom[3463] = 1;
     rom[3464] = 1;
     rom[3465] = 1;
     rom[3466] = 1;
     rom[3467] = 1;
     rom[3468] = 1;
     rom[3469] = 1;
     rom[3470] = 1;
     rom[3471] = 1;
     rom[3472] = 1;
     rom[3473] = 1;
     rom[3474] = 1;
     rom[3475] = 1;
     rom[3476] = 0;
     rom[3477] = 0;
     rom[3478] = 0;
     rom[3479] = 0;
     rom[3480] = 0;
     rom[3481] = 0;
     rom[3482] = 1;
     rom[3483] = 1;
     rom[3484] = 1;
     rom[3485] = 1;
     rom[3486] = 1;
     rom[3487] = 1;
     rom[3488] = 1;
     rom[3489] = 1;
     rom[3490] = 1;
     rom[3491] = 1;
     rom[3492] = 1;
     rom[3493] = 1;
     rom[3494] = 0;
     rom[3495] = 0;
     rom[3496] = 0;
     rom[3497] = 0;
     rom[3498] = 0;
     rom[3499] = 0;
     rom[3500] = 1;
     rom[3501] = 1;
     rom[3502] = 1;
     rom[3503] = 1;
     rom[3504] = 1;
     rom[3505] = 1;
     rom[3506] = 1;
     rom[3507] = 1;
     rom[3508] = 1;
     rom[3509] = 1;
     rom[3510] = 1;
     rom[3511] = 1;
     rom[3512] = 1;
     rom[3513] = 0;
     rom[3514] = 0;
     rom[3515] = 0;
     rom[3516] = 0;
     rom[3517] = 0;
     rom[3518] = 0;
     rom[3519] = 0;
     rom[3520] = 0;
     rom[3521] = 0;
     rom[3522] = 0;
     rom[3523] = 0;
     rom[3524] = 0;
     rom[3525] = 0;
     rom[3526] = 0;
     rom[3527] = 0;
     rom[3528] = 1;
     rom[3529] = 1;
     rom[3530] = 1;
     rom[3531] = 1;
     rom[3532] = 1;
     rom[3533] = 1;
     rom[3534] = 1;
     rom[3535] = 1;
     rom[3536] = 1;
     rom[3537] = 1;
     rom[3538] = 1;
     rom[3539] = 0;
     rom[3540] = 0;
     rom[3541] = 0;
     rom[3542] = 0;
     rom[3543] = 0;
     rom[3544] = 0;
     rom[3545] = 0;
     rom[3546] = 1;
     rom[3547] = 1;
     rom[3548] = 1;
     rom[3549] = 1;
     rom[3550] = 1;
     rom[3551] = 1;
     rom[3552] = 1;
     rom[3553] = 1;
     rom[3554] = 1;
     rom[3555] = 1;
     rom[3556] = 1;
     rom[3557] = 0;
     rom[3558] = 0;
     rom[3559] = 0;
     rom[3560] = 0;
     rom[3561] = 0;
     rom[3562] = 0;
     rom[3563] = 0;
     rom[3564] = 0;
     rom[3565] = 1;
     rom[3566] = 1;
     rom[3567] = 1;
     rom[3568] = 1;
     rom[3569] = 1;
     rom[3570] = 1;
     rom[3571] = 1;
     rom[3572] = 1;
     rom[3573] = 1;
     rom[3574] = 1;
     rom[3575] = 1;
     rom[3576] = 0;
     rom[3577] = 0;
     rom[3578] = 0;
     rom[3579] = 0;
     rom[3580] = 0;
     rom[3581] = 0;
     rom[3582] = 0;
     rom[3583] = 0;
     rom[3584] = 0;
     rom[3585] = 0;
     rom[3586] = 0;
     rom[3587] = 0;
     rom[3588] = 0;
     rom[3589] = 0;
     rom[3590] = 0;
     rom[3591] = 0;
     rom[3592] = 0;
     rom[3593] = 1;
     rom[3594] = 1;
     rom[3595] = 1;
     rom[3596] = 1;
     rom[3597] = 1;
     rom[3598] = 1;
     rom[3599] = 1;
     rom[3600] = 1;
     rom[3601] = 1;
     rom[3602] = 0;
     rom[3603] = 0;
     rom[3604] = 0;
     rom[3605] = 0;
     rom[3606] = 0;
     rom[3607] = 0;
     rom[3608] = 0;
     rom[3609] = 0;
     rom[3610] = 0;
     rom[3611] = 1;
     rom[3612] = 1;
     rom[3613] = 1;
     rom[3614] = 1;
     rom[3615] = 1;
     rom[3616] = 1;
     rom[3617] = 1;
     rom[3618] = 1;
     rom[3619] = 1;
     rom[3620] = 0;
     rom[3621] = 0;
     rom[3622] = 0;
     rom[3623] = 0;
     rom[3624] = 0;
     rom[3625] = 0;
     rom[3626] = 0;
     rom[3627] = 0;
     rom[3628] = 0;
     rom[3629] = 0;
     rom[3630] = 1;
     rom[3631] = 1;
     rom[3632] = 1;
     rom[3633] = 1;
     rom[3634] = 1;
     rom[3635] = 1;
     rom[3636] = 1;
     rom[3637] = 1;
     rom[3638] = 1;
     rom[3639] = 0;
     rom[3640] = 0;
     rom[3641] = 0;
     rom[3642] = 0;
     rom[3643] = 0;
     rom[3644] = 0;
     rom[3645] = 0;
     rom[3646] = 0;
     rom[3647] = 0;
     rom[3648] = 0;
     rom[3649] = 0;
     rom[3650] = 0;
     rom[3651] = 0;
     rom[3652] = 0;
     rom[3653] = 0;
     rom[3654] = 0;
     rom[3655] = 0;
     rom[3656] = 0;
     rom[3657] = 0;
     rom[3658] = 0;
     rom[3659] = 1;
     rom[3660] = 1;
     rom[3661] = 1;
     rom[3662] = 1;
     rom[3663] = 1;
     rom[3664] = 0;
     rom[3665] = 0;
     rom[3666] = 0;
     rom[3667] = 0;
     rom[3668] = 0;
     rom[3669] = 0;
     rom[3670] = 0;
     rom[3671] = 0;
     rom[3672] = 0;
     rom[3673] = 0;
     rom[3674] = 0;
     rom[3675] = 0;
     rom[3676] = 0;
     rom[3677] = 1;
     rom[3678] = 1;
     rom[3679] = 1;
     rom[3680] = 1;
     rom[3681] = 1;
     rom[3682] = 1;
     rom[3683] = 0;
     rom[3684] = 0;
     rom[3685] = 0;
     rom[3686] = 0;
     rom[3687] = 0;
     rom[3688] = 0;
     rom[3689] = 0;
     rom[3690] = 0;
     rom[3691] = 0;
     rom[3692] = 0;
     rom[3693] = 0;
     rom[3694] = 0;
     rom[3695] = 0;
     rom[3696] = 1;
     rom[3697] = 1;
     rom[3698] = 1;
     rom[3699] = 1;
     rom[3700] = 1;
     rom[3701] = 0;
     rom[3702] = 0;
     rom[3703] = 0;
     rom[3704] = 0;
     rom[3705] = 0;
     rom[3706] = 0;
     rom[3707] = 0;
     rom[3708] = 0;
     rom[3709] = 0;
     rom[3710] = 0;
     rom[3711] = 0;
     rom[3712] = 0;
     rom[3713] = 0;
     rom[3714] = 0;
     rom[3715] = 0;
     rom[3716] = 0;
     rom[3717] = 0;
     rom[3718] = 0;
     rom[3719] = 0;
     rom[3720] = 0;
     rom[3721] = 0;
     rom[3722] = 0;
     rom[3723] = 0;
     rom[3724] = 0;
     rom[3725] = 0;
     rom[3726] = 0;
     rom[3727] = 0;
     rom[3728] = 0;
     rom[3729] = 0;
     rom[3730] = 0;
     rom[3731] = 0;
     rom[3732] = 0;
     rom[3733] = 0;
     rom[3734] = 0;
     rom[3735] = 0;
     rom[3736] = 0;
     rom[3737] = 0;
     rom[3738] = 0;
     rom[3739] = 0;
     rom[3740] = 0;
     rom[3741] = 0;
     rom[3742] = 0;
     rom[3743] = 0;
     rom[3744] = 0;
     rom[3745] = 0;
     rom[3746] = 0;
     rom[3747] = 0;
     rom[3748] = 0;
     rom[3749] = 0;
     rom[3750] = 0;
     rom[3751] = 0;
     rom[3752] = 0;
     rom[3753] = 0;
     rom[3754] = 0;
     rom[3755] = 0;
     rom[3756] = 0;
     rom[3757] = 0;
     rom[3758] = 0;
     rom[3759] = 0;
     rom[3760] = 0;
     rom[3761] = 0;
     rom[3762] = 0;
     rom[3763] = 0;
     rom[3764] = 0;
     rom[3765] = 0;
     rom[3766] = 0;
     rom[3767] = 0;
     rom[3768] = 0;
     rom[3769] = 0;
     rom[3770] = 0;
     rom[3771] = 0;
     rom[3772] = 0;
     rom[3773] = 0;
     rom[3774] = 0;
     rom[3775] = 0;
     rom[3776] = 0;
     rom[3777] = 0;
     rom[3778] = 0;
     rom[3779] = 0;
     rom[3780] = 0;
     rom[3781] = 0;
     rom[3782] = 0;
     rom[3783] = 0;
     rom[3784] = 0;
     rom[3785] = 0;
     rom[3786] = 0;
     rom[3787] = 0;
     rom[3788] = 0;
     rom[3789] = 0;
     rom[3790] = 0;
     rom[3791] = 0;
     rom[3792] = 0;
     rom[3793] = 0;
     rom[3794] = 0;
     rom[3795] = 0;
     rom[3796] = 0;
     rom[3797] = 0;
     rom[3798] = 0;
     rom[3799] = 0;
     rom[3800] = 0;
     rom[3801] = 0;
     rom[3802] = 0;
     rom[3803] = 0;
     rom[3804] = 0;
     rom[3805] = 0;
     rom[3806] = 0;
     rom[3807] = 0;
     rom[3808] = 0;
     rom[3809] = 0;
     rom[3810] = 0;
     rom[3811] = 0;
     rom[3812] = 0;
     rom[3813] = 0;
     rom[3814] = 0;
     rom[3815] = 0;
     rom[3816] = 0;
     rom[3817] = 0;
     rom[3818] = 0;
     rom[3819] = 0;
     rom[3820] = 0;
     rom[3821] = 0;
     rom[3822] = 0;
     rom[3823] = 0;
     rom[3824] = 0;
     rom[3825] = 0;
     rom[3826] = 0;
     rom[3827] = 0;
     rom[3828] = 0;
     rom[3829] = 0;
     rom[3830] = 0;
     rom[3831] = 0;
     rom[3832] = 0;
     rom[3833] = 0;
     rom[3834] = 0;
     rom[3835] = 0;
     rom[3836] = 0;
     rom[3837] = 0;
     rom[3838] = 0;
     rom[3839] = 0;
     rom[3840] = 0;
     rom[3841] = 0;
     rom[3842] = 0;
     rom[3843] = 0;
     rom[3844] = 0;
     rom[3845] = 0;
     rom[3846] = 0;
     rom[3847] = 0;
     rom[3848] = 0;
     rom[3849] = 0;
     rom[3850] = 0;
     rom[3851] = 0;
     rom[3852] = 0;
     rom[3853] = 0;
     rom[3854] = 0;
     rom[3855] = 0;
     rom[3856] = 0;
     rom[3857] = 0;
     rom[3858] = 0;
     rom[3859] = 0;
     rom[3860] = 0;
     rom[3861] = 0;
     rom[3862] = 0;
     rom[3863] = 0;
     rom[3864] = 0;
     rom[3865] = 0;
     rom[3866] = 0;
     rom[3867] = 0;
     rom[3868] = 0;
     rom[3869] = 0;
     rom[3870] = 0;
     rom[3871] = 0;
     rom[3872] = 0;
     rom[3873] = 0;
     rom[3874] = 0;
     rom[3875] = 0;
     rom[3876] = 0;
     rom[3877] = 0;
     rom[3878] = 0;
     rom[3879] = 0;
     rom[3880] = 0;
     rom[3881] = 0;
     rom[3882] = 0;
     rom[3883] = 0;
     rom[3884] = 0;
     rom[3885] = 0;
     rom[3886] = 0;
     rom[3887] = 0;
     rom[3888] = 0;
     rom[3889] = 0;
     rom[3890] = 0;
     rom[3891] = 0;
     rom[3892] = 0;
     rom[3893] = 0;
     rom[3894] = 0;
     rom[3895] = 0;
     rom[3896] = 0;
     rom[3897] = 0;
     rom[3898] = 0;
     rom[3899] = 0;
     rom[3900] = 0;
     rom[3901] = 0;
     rom[3902] = 0;
     rom[3903] = 0;
     rom[3904] = 0;
     rom[3905] = 0;
     rom[3906] = 0;
     rom[3907] = 0;
     rom[3908] = 0;
     rom[3909] = 0;
     rom[3910] = 0;
     rom[3911] = 0;
     rom[3912] = 0;
     rom[3913] = 0;
     rom[3914] = 0;
     rom[3915] = 0;
     rom[3916] = 0;
     rom[3917] = 0;
     rom[3918] = 0;
     rom[3919] = 0;
     rom[3920] = 0;
     rom[3921] = 0;
     rom[3922] = 0;
     rom[3923] = 0;
     rom[3924] = 0;
     rom[3925] = 0;
     rom[3926] = 0;
     rom[3927] = 0;
     rom[3928] = 0;
     rom[3929] = 0;
     rom[3930] = 0;
     rom[3931] = 0;
     rom[3932] = 0;
     rom[3933] = 0;
     rom[3934] = 0;
     rom[3935] = 0;
     rom[3936] = 0;
     rom[3937] = 0;
     rom[3938] = 0;
     rom[3939] = 0;
     rom[3940] = 0;
     rom[3941] = 0;
     rom[3942] = 0;
     rom[3943] = 0;
     rom[3944] = 0;
     rom[3945] = 0;
     rom[3946] = 0;
     rom[3947] = 0;
     rom[3948] = 0;
     rom[3949] = 0;
     rom[3950] = 0;
     rom[3951] = 0;
     rom[3952] = 0;
     rom[3953] = 0;
     rom[3954] = 0;
     rom[3955] = 0;
     rom[3956] = 0;
     rom[3957] = 0;
     rom[3958] = 0;
     rom[3959] = 0;
     rom[3960] = 0;
     rom[3961] = 0;
     rom[3962] = 0;
     rom[3963] = 0;
     rom[3964] = 0;
     rom[3965] = 0;
     rom[3966] = 0;
     rom[3967] = 0;
     rom[3968] = 0;
     rom[3969] = 0;
     rom[3970] = 0;
     rom[3971] = 0;
     rom[3972] = 0;
     rom[3973] = 0;
     rom[3974] = 0;
     rom[3975] = 0;
     rom[3976] = 0;
     rom[3977] = 0;
     rom[3978] = 0;
     rom[3979] = 0;
     rom[3980] = 0;
     rom[3981] = 0;
     rom[3982] = 0;
     rom[3983] = 0;
     rom[3984] = 0;
     rom[3985] = 0;
     rom[3986] = 0;
     rom[3987] = 0;
     rom[3988] = 0;
     rom[3989] = 0;
     rom[3990] = 0;
     rom[3991] = 0;
     rom[3992] = 0;
     rom[3993] = 0;
     rom[3994] = 0;
     rom[3995] = 0;
     rom[3996] = 0;
     rom[3997] = 0;
     rom[3998] = 0;
     rom[3999] = 0;
     rom[4000] = 0;
     rom[4001] = 0;
     rom[4002] = 0;
     rom[4003] = 0;
     rom[4004] = 0;
     rom[4005] = 0;
     rom[4006] = 0;
     rom[4007] = 0;
     rom[4008] = 0;
     rom[4009] = 0;
     rom[4010] = 0;
     rom[4011] = 0;
     rom[4012] = 0;
     rom[4013] = 0;
     rom[4014] = 0;
     rom[4015] = 0;
     rom[4016] = 0;
     rom[4017] = 0;
     rom[4018] = 0;
     rom[4019] = 0;
     rom[4020] = 0;
     rom[4021] = 0;
     rom[4022] = 0;
     rom[4023] = 0;
     rom[4024] = 0;
     rom[4025] = 0;
     rom[4026] = 0;
     rom[4027] = 0;
     rom[4028] = 0;
     rom[4029] = 0;
     rom[4030] = 0;
     rom[4031] = 0;
     rom[4032] = 0;
     rom[4033] = 0;
     rom[4034] = 0;
     rom[4035] = 0;
     rom[4036] = 0;
     rom[4037] = 0;
     rom[4038] = 0;
     rom[4039] = 0;
     rom[4040] = 0;
     rom[4041] = 0;
     rom[4042] = 0;
     rom[4043] = 0;
     rom[4044] = 0;
     rom[4045] = 0;
     rom[4046] = 0;
     rom[4047] = 0;
     rom[4048] = 0;
     rom[4049] = 0;
     rom[4050] = 0;
     rom[4051] = 0;
     rom[4052] = 0;
     rom[4053] = 0;
     rom[4054] = 0;
     rom[4055] = 0;
     rom[4056] = 0;
     rom[4057] = 0;
     rom[4058] = 0;
     rom[4059] = 0;
     rom[4060] = 0;
     rom[4061] = 0;
     rom[4062] = 0;
     rom[4063] = 0;
     rom[4064] = 0;
     rom[4065] = 0;
     rom[4066] = 0;
     rom[4067] = 0;
     rom[4068] = 0;
     rom[4069] = 0;
     rom[4070] = 0;
     rom[4071] = 0;
     rom[4072] = 0;
     rom[4073] = 0;
     rom[4074] = 0;
     rom[4075] = 0;
     rom[4076] = 0;
     rom[4077] = 0;
     rom[4078] = 0;
     rom[4079] = 0;
     rom[4080] = 0;
     rom[4081] = 0;
     rom[4082] = 0;
     rom[4083] = 0;
     rom[4084] = 0;
     rom[4085] = 0;
     rom[4086] = 0;
     rom[4087] = 0;
     rom[4088] = 0;
     rom[4089] = 0;
     rom[4090] = 0;
     rom[4091] = 0;
     rom[4092] = 0;
     rom[4093] = 0;
     rom[4094] = 0;
     rom[4095] = 0;

	end

	always @ (posedge clk)
	begin
		q <= rom[addr];
	end

endmodule
